Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity violin_lut is
    generic (
        DEPTH : integer := 2048;
        WIDTH : integer := 16
    );
    port (
        clk   : in  std_logic;
        addr  : in  std_logic_vector(10 downto 0);
        dout  : out std_logic_vector(WIDTH-1 downto 0)
    );
end violin_lut;

architecture arch of violin_lut is
    type lut_array is array(0 to DEPTH-1) of std_logic_vector(WIDTH-1 downto 0);
    signal lut: lut_array := (
x"0000",
x"01D3",
x"03A7",
x"057A",
x"074D",
x"0920",
x"0AF2",
x"0CC4",
x"0E95",
x"1065",
x"1234",
x"1402",
x"15CF",
x"179B",
x"1966",
x"1B2F",
x"1CF7",
x"1EBD",
x"2082",
x"2245",
x"2406",
x"25C5",
x"2782",
x"293D",
x"2AF5",
x"2CAC",
x"2E60",
x"3012",
x"31C1",
x"336D",
x"3517",
x"36BE",
x"3862",
x"3A03",
x"3BA1",
x"3D3C",
x"3ED4",
x"4068",
x"41F9",
x"4387",
x"4512",
x"4699",
x"481C",
x"499B",
x"4B17",
x"4C90",
x"4E04",
x"4F74",
x"50E1",
x"5249",
x"53AE",
x"550E",
x"566A",
x"57C2",
x"5916",
x"5A65",
x"5BB1",
x"5CF7",
x"5E3A",
x"5F78",
x"60B1",
x"61E6",
x"6317",
x"6442",
x"656A",
x"668C",
x"67AB",
x"68C4",
x"69D9",
x"6AE9",
x"6BF4",
x"6CFB",
x"6DFD",
x"6EFA",
x"6FF2",
x"70E6",
x"71D5",
x"72BF",
x"73A5",
x"7485",
x"7561",
x"7638",
x"770B",
x"77D9",
x"78A2",
x"7966",
x"7A25",
x"7AE0",
x"7B97",
x"7C48",
x"7CF5",
x"7D9E",
x"7E42",
x"7EE1",
x"7F7C",
x"8012",
x"80A4",
x"8131",
x"81BA",
x"823F",
x"82BF",
x"833B",
x"83B3",
x"8427",
x"8496",
x"8501",
x"8568",
x"85CB",
x"862B",
x"8686",
x"86DD",
x"8730",
x"8780",
x"87CC",
x"8814",
x"8858",
x"8899",
x"88D7",
x"8911",
x"8947",
x"897A",
x"89AA",
x"89D6",
x"89FF",
x"8A25",
x"8A48",
x"8A68",
x"8A85",
x"8A9F",
x"8AB7",
x"8ACB",
x"8ADD",
x"8AEC",
x"8AF8",
x"8B02",
x"8B09",
x"8B0E",
x"8B11",
x"8B11",
x"8B0F",
x"8B0B",
x"8B05",
x"8AFD",
x"8AF3",
x"8AE6",
x"8AD8",
x"8AC9",
x"8AB7",
x"8AA4",
x"8A8F",
x"8A78",
x"8A60",
x"8A47",
x"8A2C",
x"8A10",
x"89F3",
x"89D4",
x"89B5",
x"8994",
x"8972",
x"894F",
x"892B",
x"8907",
x"88E1",
x"88BB",
x"8894",
x"886D",
x"8844",
x"881C",
x"87F2",
x"87C8",
x"879E",
x"8774",
x"8749",
x"871D",
x"86F2",
x"86C6",
x"869A",
x"866F",
x"8642",
x"8616",
x"85EA",
x"85BE",
x"8592",
x"8566",
x"853A",
x"850F",
x"84E3",
x"84B8",
x"848D",
x"8463",
x"8438",
x"840E",
x"83E5",
x"83BB",
x"8393",
x"836A",
x"8342",
x"831B",
x"82F4",
x"82CD",
x"82A7",
x"8282",
x"825D",
x"8239",
x"8215",
x"81F2",
x"81D0",
x"81AE",
x"818D",
x"816D",
x"814D",
x"812E",
x"810F",
x"80F1",
x"80D4",
x"80B8",
x"809C",
x"8081",
x"8066",
x"804C",
x"8033",
x"801B",
x"8003",
x"7FEC",
x"7FD6",
x"7FC0",
x"7FAB",
x"7F97",
x"7F84",
x"7F71",
x"7F5E",
x"7F4D",
x"7F3B",
x"7F2B",
x"7F1B",
x"7F0C",
x"7EFD",
x"7EEF",
x"7EE2",
x"7ED5",
x"7EC8",
x"7EBD",
x"7EB1",
x"7EA7",
x"7E9C",
x"7E92",
x"7E89",
x"7E80",
x"7E78",
x"7E70",
x"7E68",
x"7E61",
x"7E5A",
x"7E54",
x"7E4E",
x"7E48",
x"7E42",
x"7E3D",
x"7E38",
x"7E34",
x"7E30",
x"7E2C",
x"7E28",
x"7E24",
x"7E21",
x"7E1E",
x"7E1B",
x"7E18",
x"7E15",
x"7E12",
x"7E10",
x"7E0D",
x"7E0B",
x"7E09",
x"7E07",
x"7E04",
x"7E02",
x"7E00",
x"7DFE",
x"7DFC",
x"7DFA",
x"7DF7",
x"7DF5",
x"7DF3",
x"7DF0",
x"7DEE",
x"7DEB",
x"7DE8",
x"7DE6",
x"7DE3",
x"7DE0",
x"7DDC",
x"7DD9",
x"7DD5",
x"7DD2",
x"7DCE",
x"7DCA",
x"7DC5",
x"7DC1",
x"7DBC",
x"7DB7",
x"7DB2",
x"7DAD",
x"7DA7",
x"7DA1",
x"7D9B",
x"7D95",
x"7D8E",
x"7D87",
x"7D80",
x"7D79",
x"7D72",
x"7D6A",
x"7D62",
x"7D59",
x"7D51",
x"7D48",
x"7D3F",
x"7D35",
x"7D2C",
x"7D22",
x"7D18",
x"7D0D",
x"7D02",
x"7CF8",
x"7CEC",
x"7CE1",
x"7CD5",
x"7CC9",
x"7CBD",
x"7CB1",
x"7CA4",
x"7C97",
x"7C8A",
x"7C7D",
x"7C70",
x"7C62",
x"7C54",
x"7C46",
x"7C38",
x"7C29",
x"7C1B",
x"7C0C",
x"7BFD",
x"7BEE",
x"7BDE",
x"7BCF",
x"7BBF",
x"7BB0",
x"7BA0",
x"7B90",
x"7B80",
x"7B6F",
x"7B5F",
x"7B4F",
x"7B3E",
x"7B2D",
x"7B1D",
x"7B0C",
x"7AFB",
x"7AEA",
x"7AD9",
x"7AC8",
x"7AB7",
x"7AA6",
x"7A95",
x"7A84",
x"7A73",
x"7A62",
x"7A51",
x"7A3F",
x"7A2E",
x"7A1D",
x"7A0C",
x"79FB",
x"79EA",
x"79D9",
x"79C8",
x"79B7",
x"79A6",
x"7995",
x"7984",
x"7973",
x"7962",
x"7951",
x"7941",
x"7930",
x"7920",
x"790F",
x"78FF",
x"78EE",
x"78DE",
x"78CE",
x"78BE",
x"78AE",
x"789E",
x"788E",
x"787E",
x"786E",
x"785F",
x"784F",
x"783F",
x"7830",
x"7820",
x"7811",
x"7802",
x"77F3",
x"77E3",
x"77D4",
x"77C5",
x"77B6",
x"77A7",
x"7798",
x"7789",
x"777B",
x"776C",
x"775D",
x"774E",
x"7740",
x"7731",
x"7722",
x"7714",
x"7705",
x"76F6",
x"76E7",
x"76D9",
x"76CA",
x"76BB",
x"76AD",
x"769E",
x"768F",
x"7680",
x"7671",
x"7662",
x"7653",
x"7644",
x"7635",
x"7625",
x"7616",
x"7606",
x"75F7",
x"75E7",
x"75D7",
x"75C7",
x"75B7",
x"75A7",
x"7597",
x"7586",
x"7575",
x"7565",
x"7554",
x"7542",
x"7531",
x"751F",
x"750E",
x"74FC",
x"74E9",
x"74D7",
x"74C5",
x"74B2",
x"749F",
x"748B",
x"7478",
x"7464",
x"7450",
x"743C",
x"7427",
x"7412",
x"73FD",
x"73E8",
x"73D2",
x"73BC",
x"73A6",
x"7390",
x"7379",
x"7362",
x"734A",
x"7333",
x"731B",
x"7302",
x"72EA",
x"72D1",
x"72B8",
x"729E",
x"7284",
x"726A",
x"724F",
x"7235",
x"7219",
x"71FE",
x"71E2",
x"71C6",
x"71AA",
x"718D",
x"7170",
x"7153",
x"7135",
x"7117",
x"70F8",
x"70DA",
x"70BB",
x"709C",
x"707C",
x"705C",
x"703C",
x"701C",
x"6FFB",
x"6FDA",
x"6FB9",
x"6F97",
x"6F75",
x"6F53",
x"6F31",
x"6F0E",
x"6EEB",
x"6EC8",
x"6EA5",
x"6E81",
x"6E5D",
x"6E39",
x"6E14",
x"6DF0",
x"6DCB",
x"6DA6",
x"6D81",
x"6D5C",
x"6D36",
x"6D10",
x"6CEA",
x"6CC4",
x"6C9E",
x"6C77",
x"6C51",
x"6C2A",
x"6C03",
x"6BDC",
x"6BB5",
x"6B8E",
x"6B66",
x"6B3F",
x"6B17",
x"6AF0",
x"6AC8",
x"6AA0",
x"6A78",
x"6A51",
x"6A29",
x"6A01",
x"69D8",
x"69B0",
x"6988",
x"6960",
x"6938",
x"6910",
x"68E8",
x"68C0",
x"6897",
x"686F",
x"6847",
x"681F",
x"67F7",
x"67CF",
x"67A7",
x"677F",
x"6758",
x"6730",
x"6708",
x"66E1",
x"66B9",
x"6692",
x"666A",
x"6643",
x"661C",
x"65F5",
x"65CE",
x"65A7",
x"6580",
x"6559",
x"6533",
x"650D",
x"64E6",
x"64C0",
x"649A",
x"6474",
x"644E",
x"6429",
x"6403",
x"63DE",
x"63B8",
x"6393",
x"636E",
x"6349",
x"6324",
x"6300",
x"62DB",
x"62B7",
x"6293",
x"626F",
x"624B",
x"6227",
x"6203",
x"61DF",
x"61BC",
x"6198",
x"6175",
x"6152",
x"612F",
x"610C",
x"60E9",
x"60C6",
x"60A3",
x"6081",
x"605E",
x"603C",
x"601A",
x"5FF7",
x"5FD5",
x"5FB3",
x"5F91",
x"5F6F",
x"5F4D",
x"5F2B",
x"5F09",
x"5EE7",
x"5EC5",
x"5EA3",
x"5E81",
x"5E5F",
x"5E3E",
x"5E1C",
x"5DFA",
x"5DD8",
x"5DB6",
x"5D94",
x"5D72",
x"5D50",
x"5D2E",
x"5D0B",
x"5CE9",
x"5CC7",
x"5CA4",
x"5C82",
x"5C5F",
x"5C3D",
x"5C1A",
x"5BF7",
x"5BD4",
x"5BB0",
x"5B8D",
x"5B6A",
x"5B46",
x"5B22",
x"5AFE",
x"5ADA",
x"5AB6",
x"5A91",
x"5A6C",
x"5A47",
x"5A22",
x"59FD",
x"59D7",
x"59B1",
x"598B",
x"5965",
x"593F",
x"5918",
x"58F1",
x"58C9",
x"58A2",
x"587A",
x"5852",
x"5829",
x"5801",
x"57D8",
x"57AF",
x"5785",
x"575B",
x"5731",
x"5706",
x"56DB",
x"56B0",
x"5685",
x"5659",
x"562D",
x"5600",
x"55D4",
x"55A6",
x"5579",
x"554B",
x"551D",
x"54EE",
x"54C0",
x"5490",
x"5461",
x"5431",
x"5401",
x"53D0",
x"539F",
x"536E",
x"533C",
x"530A",
x"52D7",
x"52A5",
x"5272",
x"523E",
x"520A",
x"51D6",
x"51A2",
x"516D",
x"5137",
x"5102",
x"50CC",
x"5096",
x"505F",
x"5028",
x"4FF1",
x"4FB9",
x"4F81",
x"4F49",
x"4F11",
x"4ED8",
x"4E9F",
x"4E65",
x"4E2B",
x"4DF1",
x"4DB7",
x"4D7C",
x"4D41",
x"4D06",
x"4CCA",
x"4C8E",
x"4C52",
x"4C16",
x"4BD9",
x"4B9C",
x"4B5F",
x"4B21",
x"4AE4",
x"4AA6",
x"4A67",
x"4A29",
x"49EA",
x"49AB",
x"496C",
x"492D",
x"48EE",
x"48AE",
x"486E",
x"482E",
x"47ED",
x"47AD",
x"476C",
x"472C",
x"46EB",
x"46A9",
x"4668",
x"4627",
x"45E5",
x"45A3",
x"4561",
x"451F",
x"44DD",
x"449B",
x"4459",
x"4416",
x"43D4",
x"4391",
x"434E",
x"430B",
x"42C8",
x"4285",
x"4242",
x"41FF",
x"41BC",
x"4178",
x"4135",
x"40F2",
x"40AE",
x"406A",
x"4027",
x"3FE3",
x"3F9F",
x"3F5C",
x"3F18",
x"3ED4",
x"3E90",
x"3E4C",
x"3E09",
x"3DC5",
x"3D81",
x"3D3D",
x"3CF9",
x"3CB5",
x"3C71",
x"3C2D",
x"3BE9",
x"3BA5",
x"3B61",
x"3B1D",
x"3AD9",
x"3A95",
x"3A51",
x"3A0D",
x"39C9",
x"3985",
x"3941",
x"38FD",
x"38B9",
x"3875",
x"3831",
x"37ED",
x"37A9",
x"3765",
x"3721",
x"36DD",
x"3699",
x"3655",
x"3611",
x"35CD",
x"3589",
x"3545",
x"3502",
x"34BE",
x"347A",
x"3436",
x"33F2",
x"33AE",
x"336A",
x"3326",
x"32E2",
x"329E",
x"325B",
x"3217",
x"31D3",
x"318F",
x"314B",
x"3107",
x"30C3",
x"307F",
x"303B",
x"2FF7",
x"2FB3",
x"2F6F",
x"2F2A",
x"2EE6",
x"2EA2",
x"2E5E",
x"2E1A",
x"2DD6",
x"2D91",
x"2D4D",
x"2D09",
x"2CC4",
x"2C80",
x"2C3B",
x"2BF7",
x"2BB2",
x"2B6E",
x"2B29",
x"2AE5",
x"2AA0",
x"2A5B",
x"2A16",
x"29D2",
x"298D",
x"2948",
x"2903",
x"28BE",
x"2879",
x"2834",
x"27EF",
x"27A9",
x"2764",
x"271F",
x"26D9",
x"2694",
x"264F",
x"2609",
x"25C4",
x"257E",
x"2538",
x"24F3",
x"24AD",
x"2467",
x"2421",
x"23DB",
x"2395",
x"2350",
x"230A",
x"22C4",
x"227D",
x"2237",
x"21F1",
x"21AB",
x"2165",
x"211F",
x"20D8",
x"2092",
x"204C",
x"2005",
x"1FBF",
x"1F79",
x"1F32",
x"1EEC",
x"1EA5",
x"1E5F",
x"1E18",
x"1DD2",
x"1D8C",
x"1D45",
x"1CFF",
x"1CB8",
x"1C72",
x"1C2B",
x"1BE5",
x"1B9F",
x"1B58",
x"1B12",
x"1ACC",
x"1A85",
x"1A3F",
x"19F9",
x"19B2",
x"196C",
x"1926",
x"18E0",
x"189A",
x"1854",
x"180E",
x"17C8",
x"1782",
x"173D",
x"16F7",
x"16B1",
x"166C",
x"1626",
x"15E1",
x"159C",
x"1556",
x"1511",
x"14CC",
x"1487",
x"1442",
x"13FD",
x"13B9",
x"1374",
x"1330",
x"12EB",
x"12A7",
x"1263",
x"121F",
x"11DB",
x"1197",
x"1153",
x"110F",
x"10CC",
x"1088",
x"1045",
x"1002",
x"0FBF",
x"0F7C",
x"0F39",
x"0EF6",
x"0EB4",
x"0E71",
x"0E2F",
x"0DED",
x"0DAB",
x"0D69",
x"0D27",
x"0CE6",
x"0CA4",
x"0C63",
x"0C21",
x"0BE0",
x"0B9F",
x"0B5E",
x"0B1D",
x"0ADD",
x"0A9C",
x"0A5C",
x"0A1C",
x"09DB",
x"099B",
x"095B",
x"091C",
x"08DC",
x"089C",
x"085D",
x"081D",
x"07DE",
x"079F",
x"0760",
x"0721",
x"06E2",
x"06A3",
x"0665",
x"0626",
x"05E8",
x"05A9",
x"056B",
x"052D",
x"04EF",
x"04B1",
x"0472",
x"0435",
x"03F7",
x"03B9",
x"037B",
x"033D",
x"0300",
x"02C2",
x"0284",
x"0247",
x"0209",
x"01CC",
x"018E",
x"0151",
x"0114",
x"00D6",
x"0099",
x"005C",
x"001E",
x"FFE2",
x"FFA4",
x"FF67",
x"FF2A",
x"FEEC",
x"FEAF",
x"FE72",
x"FE34",
x"FDF7",
x"FDB9",
x"FD7C",
x"FD3E",
x"FD00",
x"FCC3",
x"FC85",
x"FC47",
x"FC09",
x"FBCB",
x"FB8E",
x"FB4F",
x"FB11",
x"FAD3",
x"FA95",
x"FA57",
x"FA18",
x"F9DA",
x"F99B",
x"F95D",
x"F91E",
x"F8DF",
x"F8A0",
x"F861",
x"F822",
x"F7E3",
x"F7A3",
x"F764",
x"F724",
x"F6E4",
x"F6A5",
x"F665",
x"F625",
x"F5E4",
x"F5A4",
x"F564",
x"F523",
x"F4E3",
x"F4A2",
x"F461",
x"F420",
x"F3DF",
x"F39D",
x"F35C",
x"F31A",
x"F2D9",
x"F297",
x"F255",
x"F213",
x"F1D1",
x"F18F",
x"F14C",
x"F10A",
x"F0C7",
x"F084",
x"F041",
x"EFFE",
x"EFBB",
x"EF78",
x"EF34",
x"EEF1",
x"EEAD",
x"EE69",
x"EE25",
x"EDE1",
x"ED9D",
x"ED59",
x"ED15",
x"ECD0",
x"EC8C",
x"EC47",
x"EC03",
x"EBBE",
x"EB79",
x"EB34",
x"EAEF",
x"EAAA",
x"EA64",
x"EA1F",
x"E9DA",
x"E994",
x"E94F",
x"E909",
x"E8C3",
x"E87E",
x"E838",
x"E7F2",
x"E7AC",
x"E766",
x"E720",
x"E6DA",
x"E694",
x"E64E",
x"E607",
x"E5C1",
x"E57B",
x"E534",
x"E4EE",
x"E4A8",
x"E461",
x"E41B",
x"E3D5",
x"E38E",
x"E348",
x"E301",
x"E2BB",
x"E274",
x"E22E",
x"E1E8",
x"E1A1",
x"E15B",
x"E114",
x"E0CE",
x"E087",
x"E041",
x"DFFB",
x"DFB4",
x"DF6E",
x"DF28",
x"DEE1",
x"DE9B",
x"DE55",
x"DE0F",
x"DDC9",
x"DD83",
x"DD3C",
x"DCF6",
x"DCB0",
x"DC6B",
x"DC25",
x"DBDF",
x"DB99",
x"DB53",
x"DB0D",
x"DAC8",
x"DA82",
x"DA3C",
x"D9F7",
x"D9B1",
x"D96C",
x"D927",
x"D8E1",
x"D89C",
x"D857",
x"D811",
x"D7CC",
x"D787",
x"D742",
x"D6FD",
x"D6B8",
x"D673",
x"D62E",
x"D5EA",
x"D5A5",
x"D560",
x"D51B",
x"D4D7",
x"D492",
x"D44E",
x"D409",
x"D3C5",
x"D380",
x"D33C",
x"D2F7",
x"D2B3",
x"D26F",
x"D22A",
x"D1E6",
x"D1A2",
x"D15E",
x"D11A",
x"D0D6",
x"D091",
x"D04D",
x"D009",
x"CFC5",
x"CF81",
x"CF3D",
x"CEF9",
x"CEB5",
x"CE71",
x"CE2D",
x"CDE9",
x"CDA5",
x"CD62",
x"CD1E",
x"CCDA",
x"CC96",
x"CC52",
x"CC0E",
x"CBCA",
x"CB86",
x"CB42",
x"CAFE",
x"CABB",
x"CA77",
x"CA33",
x"C9EF",
x"C9AB",
x"C967",
x"C923",
x"C8DF",
x"C89B",
x"C857",
x"C813",
x"C7CF",
x"C78B",
x"C747",
x"C703",
x"C6BF",
x"C67B",
x"C637",
x"C5F3",
x"C5AF",
x"C56B",
x"C527",
x"C4E3",
x"C49F",
x"C45B",
x"C417",
x"C3D3",
x"C38F",
x"C34B",
x"C307",
x"C2C3",
x"C27F",
x"C23B",
x"C1F7",
x"C1B4",
x"C170",
x"C12C",
x"C0E8",
x"C0A4",
x"C061",
x"C01D",
x"BFD9",
x"BF96",
x"BF52",
x"BF0E",
x"BECB",
x"BE88",
x"BE44",
x"BE01",
x"BDBE",
x"BD7B",
x"BD38",
x"BCF5",
x"BCB2",
x"BC6F",
x"BC2C",
x"BBEA",
x"BBA7",
x"BB65",
x"BB23",
x"BAE1",
x"BA9F",
x"BA5D",
x"BA1B",
x"B9D9",
x"B998",
x"B957",
x"B915",
x"B8D4",
x"B894",
x"B853",
x"B813",
x"B7D2",
x"B792",
x"B752",
x"B712",
x"B6D3",
x"B694",
x"B655",
x"B616",
x"B5D7",
x"B599",
x"B55A",
x"B51C",
x"B4DF",
x"B4A1",
x"B464",
x"B427",
x"B3EA",
x"B3AE",
x"B372",
x"B336",
x"B2FA",
x"B2BF",
x"B284",
x"B249",
x"B20F",
x"B1D5",
x"B19B",
x"B161",
x"B128",
x"B0EF",
x"B0B7",
x"B07F",
x"B047",
x"B00F",
x"AFD8",
x"AFA1",
x"AF6A",
x"AF34",
x"AEFE",
x"AEC9",
x"AE93",
x"AE5E",
x"AE2A",
x"ADF6",
x"ADC2",
x"AD8E",
x"AD5B",
x"AD29",
x"ACF6",
x"ACC4",
x"AC92",
x"AC61",
x"AC30",
x"ABFF",
x"ABCF",
x"AB9F",
x"AB70",
x"AB40",
x"AB12",
x"AAE3",
x"AAB5",
x"AA87",
x"AA5A",
x"AA2C",
x"AA00",
x"A9D3",
x"A9A7",
x"A97B",
x"A950",
x"A925",
x"A8FA",
x"A8CF",
x"A8A5",
x"A87B",
x"A851",
x"A828",
x"A7FF",
x"A7D7",
x"A7AE",
x"A786",
x"A75E",
x"A737",
x"A70F",
x"A6E8",
x"A6C1",
x"A69B",
x"A675",
x"A64F",
x"A629",
x"A603",
x"A5DE",
x"A5B9",
x"A594",
x"A56F",
x"A54A",
x"A526",
x"A502",
x"A4DE",
x"A4BA",
x"A496",
x"A473",
x"A450",
x"A42C",
x"A409",
x"A3E6",
x"A3C3",
x"A3A1",
x"A37E",
x"A35C",
x"A339",
x"A317",
x"A2F5",
x"A2D2",
x"A2B0",
x"A28E",
x"A26C",
x"A24A",
x"A228",
x"A206",
x"A1E4",
x"A1C2",
x"A1A1",
x"A17F",
x"A15D",
x"A13B",
x"A119",
x"A0F7",
x"A0D5",
x"A0B3",
x"A091",
x"A06F",
x"A04D",
x"A02B",
x"A009",
x"9FE6",
x"9FC4",
x"9FA2",
x"9F7F",
x"9F5D",
x"9F3A",
x"9F17",
x"9EF4",
x"9ED1",
x"9EAE",
x"9E8B",
x"9E68",
x"9E44",
x"9E21",
x"9DFD",
x"9DD9",
x"9DB5",
x"9D91",
x"9D6D",
x"9D49",
x"9D25",
x"9D00",
x"9CDC",
x"9CB7",
x"9C92",
x"9C6D",
x"9C48",
x"9C22",
x"9BFD",
x"9BD7",
x"9BB2",
x"9B8C",
x"9B66",
x"9B40",
x"9B1A",
x"9AF3",
x"9ACD",
x"9AA7",
x"9A80",
x"9A59",
x"9A32",
x"9A0B",
x"99E4",
x"99BD",
x"9996",
x"996E",
x"9947",
x"991F",
x"98F8",
x"98D0",
x"98A8",
x"9881",
x"9859",
x"9831",
x"9809",
x"97E1",
x"97B9",
x"9791",
x"9769",
x"9740",
x"9718",
x"96F0",
x"96C8",
x"96A0",
x"9678",
x"9650",
x"9628",
x"95FF",
x"95D7",
x"95AF",
x"9588",
x"9560",
x"9538",
x"9510",
x"94E9",
x"94C1",
x"949A",
x"9472",
x"944B",
x"9424",
x"93FD",
x"93D6",
x"93AF",
x"9389",
x"9362",
x"933C",
x"9316",
x"92F0",
x"92CA",
x"92A4",
x"927F",
x"925A",
x"9235",
x"9210",
x"91EC",
x"91C7",
x"91A3",
x"917F",
x"915B",
x"9138",
x"9115",
x"90F2",
x"90CF",
x"90AD",
x"908B",
x"9069",
x"9047",
x"9026",
x"9005",
x"8FE4",
x"8FC4",
x"8FA4",
x"8F84",
x"8F64",
x"8F45",
x"8F26",
x"8F08",
x"8EE9",
x"8ECB",
x"8EAD",
x"8E90",
x"8E73",
x"8E56",
x"8E3A",
x"8E1E",
x"8E02",
x"8DE7",
x"8DCB",
x"8DB1",
x"8D96",
x"8D7C",
x"8D62",
x"8D48",
x"8D2F",
x"8D16",
x"8CFE",
x"8CE5",
x"8CCD",
x"8CB6",
x"8C9E",
x"8C87",
x"8C70",
x"8C5A",
x"8C44",
x"8C2E",
x"8C18",
x"8C03",
x"8BEE",
x"8BD9",
x"8BC4",
x"8BB0",
x"8B9C",
x"8B88",
x"8B75",
x"8B61",
x"8B4E",
x"8B3B",
x"8B29",
x"8B17",
x"8B04",
x"8AF2",
x"8AE1",
x"8ACF",
x"8ABE",
x"8AAC",
x"8A9B",
x"8A8B",
x"8A7A",
x"8A69",
x"8A59",
x"8A49",
x"8A39",
x"8A29",
x"8A19",
x"8A09",
x"89FA",
x"89EA",
x"89DB",
x"89CB",
x"89BC",
x"89AD",
x"899E",
x"898F",
x"8980",
x"8971",
x"8962",
x"8953",
x"8945",
x"8936",
x"8927",
x"8919",
x"890A",
x"88FB",
x"88EC",
x"88DE",
x"88CF",
x"88C0",
x"88B2",
x"88A3",
x"8894",
x"8885",
x"8877",
x"8868",
x"8859",
x"884A",
x"883B",
x"882C",
x"881D",
x"880D",
x"87FE",
x"87EF",
x"87E0",
x"87D0",
x"87C1",
x"87B1",
x"87A1",
x"8792",
x"8782",
x"8772",
x"8762",
x"8752",
x"8742",
x"8732",
x"8722",
x"8712",
x"8701",
x"86F1",
x"86E0",
x"86D0",
x"86BF",
x"86AF",
x"869E",
x"868D",
x"867C",
x"866B",
x"865A",
x"8649",
x"8638",
x"8627",
x"8616",
x"8605",
x"85F4",
x"85E3",
x"85D2",
x"85C1",
x"85AF",
x"859E",
x"858D",
x"857C",
x"856B",
x"855A",
x"8549",
x"8538",
x"8527",
x"8516",
x"8505",
x"84F4",
x"84E3",
x"84D3",
x"84C2",
x"84B1",
x"84A1",
x"8491",
x"8480",
x"8470",
x"8460",
x"8450",
x"8441",
x"8431",
x"8422",
x"8412",
x"8403",
x"83F4",
x"83E5",
x"83D7",
x"83C8",
x"83BA",
x"83AC",
x"839E",
x"8390",
x"8383",
x"8376",
x"8369",
x"835C",
x"834F",
x"8343",
x"8337",
x"832B",
x"831F",
x"8314",
x"8308",
x"82FE",
x"82F3",
x"82E8",
x"82DE",
x"82D4",
x"82CB",
x"82C1",
x"82B8",
x"82AF",
x"82A7",
x"829E",
x"8296",
x"828E",
x"8287",
x"8280",
x"8279",
x"8272",
x"826B",
x"8265",
x"825F",
x"8259",
x"8253",
x"824E",
x"8249",
x"8244",
x"823F",
x"823B",
x"8236",
x"8232",
x"822E",
x"822B",
x"8227",
x"8224",
x"8220",
x"821D",
x"821A",
x"8218",
x"8215",
x"8212",
x"8210",
x"820D",
x"820B",
x"8209",
x"8206",
x"8204",
x"8202",
x"8200",
x"81FE",
x"81FC",
x"81F9",
x"81F7",
x"81F5",
x"81F3",
x"81F0",
x"81EE",
x"81EB",
x"81E8",
x"81E5",
x"81E2",
x"81DF",
x"81DC",
x"81D8",
x"81D4",
x"81D0",
x"81CC",
x"81C8",
x"81C3",
x"81BE",
x"81B8",
x"81B2",
x"81AC",
x"81A6",
x"819F",
x"8198",
x"8190",
x"8188",
x"8180",
x"8177",
x"816E",
x"8164",
x"8159",
x"814F",
x"8143",
x"8138",
x"812B",
x"811E",
x"8111",
x"8103",
x"80F4",
x"80E5",
x"80D5",
x"80C5",
x"80B3",
x"80A2",
x"808F",
x"807C",
x"8069",
x"8055",
x"8040",
x"802A",
x"8014",
x"7FFD",
x"7FE5",
x"7FCD",
x"7FB4",
x"7F9A",
x"7F7F",
x"7F64",
x"7F48",
x"7F2C",
x"7F0F",
x"7EF1",
x"7ED2",
x"7EB3",
x"7E93",
x"7E73",
x"7E52",
x"7E30",
x"7E0E",
x"7DEB",
x"7DC7",
x"7DA3",
x"7D7E",
x"7D59",
x"7D33",
x"7D0C",
x"7CE5",
x"7CBE",
x"7C96",
x"7C6D",
x"7C45",
x"7C1B",
x"7BF2",
x"7BC8",
x"7B9D",
x"7B73",
x"7B48",
x"7B1D",
x"7AF1",
x"7AC6",
x"7A9A",
x"7A6E",
x"7A42",
x"7A16",
x"79EA",
x"79BE",
x"7991",
x"7966",
x"793A",
x"790E",
x"78E3",
x"78B7",
x"788C",
x"7862",
x"7838",
x"780E",
x"77E4",
x"77BC",
x"7793",
x"776C",
x"7745",
x"771F",
x"76F9",
x"76D5",
x"76B1",
x"768E",
x"766C",
x"764B",
x"762C",
x"760D",
x"75F0",
x"75D4",
x"75B9",
x"75A0",
x"7588",
x"7571",
x"755C",
x"7549",
x"7537",
x"7528",
x"751A",
x"750D",
x"7503",
x"74FB",
x"74F5",
x"74F1",
x"74EF",
x"74EF",
x"74F2",
x"74F7",
x"74FE",
x"7508",
x"7514",
x"7523",
x"7535",
x"7549",
x"7561",
x"757B",
x"7598",
x"75B8",
x"75DB",
x"7601",
x"762A",
x"7656",
x"7686",
x"76B9",
x"76EF",
x"7729",
x"7767",
x"77A8",
x"77EC",
x"7834",
x"7880",
x"78D0",
x"7923",
x"797A",
x"79D5",
x"7A35",
x"7A98",
x"7AFF",
x"7B6A",
x"7BD9",
x"7C4D",
x"7CC5",
x"7D41",
x"7DC1",
x"7E46",
x"7ECF",
x"7F5C",
x"7FEE",
x"8084",
x"811F",
x"81BE",
x"8262",
x"830B",
x"83B8",
x"8469",
x"8520",
x"85DB",
x"869A",
x"875E",
x"8827",
x"88F5",
x"89C8",
x"8A9F",
x"8B7B",
x"8C5B",
x"8D41",
x"8E2B",
x"8F1A",
x"900E",
x"9106",
x"9203",
x"9305",
x"940C",
x"9517",
x"9627",
x"973C",
x"9855",
x"9974",
x"9A96",
x"9BBE",
x"9CE9",
x"9E1A",
x"9F4F",
x"A088",
x"A1C6",
x"A309",
x"A44F",
x"A59B",
x"A6EA",
x"A83E",
x"A996",
x"AAF2",
x"AC52",
x"ADB7",
x"AF1F",
x"B08C",
x"B1FC",
x"B370",
x"B4E9",
x"B665",
x"B7E4",
x"B967",
x"BAEE",
x"BC79",
x"BE07",
x"BF98",
x"C12C",
x"C2C4",
x"C45F",
x"C5FD",
x"C79E",
x"C942",
x"CAE9",
x"CC93",
x"CE3F",
x"CFEE",
x"D1A0",
x"D354",
x"D50B",
x"D6C3",
x"D87E",
x"DA3B",
x"DBFA",
x"DDBB",
x"DF7E",
x"E143",
x"E309",
x"E4D1",
x"E69A",
x"E865",
x"EA31",
x"EBFE",
x"EDCC",
x"EF9B",
x"F16B",
x"F33C",
x"F50E",
x"F6E0",
x"F8B3",
x"FA86",
x"FC59",
x"FE2D",
x"0000"




    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            dout <= lut(to_integer(unsigned(addr)));
        end if;
    end process;
end arch;
