Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity sine_lut is
    generic (
        DEPTH : integer := 2048;
        WIDTH : integer := 16
    );
    port (
        clk   : in  std_logic;
        addr  : in  std_logic_vector(10 downto 0);
        dout  : out std_logic_vector(WIDTH-1 downto 0)
    );
end sine_lut;

architecture arch of sine_lut is
    type lut_array is array(0 to DEPTH-1) of std_logic_vector(WIDTH-1 downto 0);
    signal lut: lut_array := (
        x"0000", x"0064", x"00C9", x"012D", x"0192", x"01F6", x"025B", x"02BF",
        x"0324", x"0388", x"03ED", x"0451", x"04B6", x"051A", x"057E", x"05E3",
        x"0647", x"06AC", x"0710", x"0774", x"07D9", x"083D", x"08A1", x"0906",
        x"096A", x"09CE", x"0A32", x"0A97", x"0AFB", x"0B5F", x"0BC3", x"0C27",
        x"0C8B", x"0CEF", x"0D53", x"0DB7", x"0E1B", x"0E7F", x"0EE3", x"0F47",
        x"0FAB", x"100E", x"1072", x"10D6", x"1139", x"119D", x"1200", x"1264",
        x"12C7", x"132B", x"138E", x"13F2", x"1455", x"14B8", x"151B", x"157E",
        x"15E1", x"1644", x"16A7", x"170A", x"176D", x"17D0", x"1833", x"1895",
        x"18F8", x"195B", x"19BD", x"1A20", x"1A82", x"1AE4", x"1B46", x"1BA9",
        x"1C0B", x"1C6D", x"1CCF", x"1D31", x"1D93", x"1DF4", x"1E56", x"1EB8",
        x"1F19", x"1F7B", x"1FDC", x"203D", x"209F", x"2100", x"2161", x"21C2",
        x"2223", x"2284", x"22E4", x"2345", x"23A6", x"2406", x"2467", x"24C7",
        x"2527", x"2587", x"25E7", x"2647", x"26A7", x"2707", x"2767", x"27C6",
        x"2826", x"2885", x"28E5", x"2944", x"29A3", x"2A02", x"2A61", x"2AC0",
        x"2B1E", x"2B7D", x"2BDB", x"2C3A", x"2C98", x"2CF6", x"2D54", x"2DB2",
        x"2E10", x"2E6E", x"2ECC", x"2F29", x"2F86", x"2FE4", x"3041", x"309E",
        x"30FB", x"3158", x"31B4", x"3211", x"326D", x"32CA", x"3326", x"3382",
        x"33DE", x"343A", x"3496", x"34F1", x"354D", x"35A8", x"3603", x"365E",
        x"36B9", x"3714", x"376F", x"37C9", x"3824", x"387E", x"38D8", x"3932",
        x"398C", x"39E6", x"3A3F", x"3A99", x"3AF2", x"3B4B", x"3BA4", x"3BFD",
        x"3C56", x"3CAE", x"3D07", x"3D5F", x"3DB7", x"3E0F", x"3E67", x"3EBF",
        x"3F16", x"3F6E", x"3FC5", x"401C", x"4073", x"40CA", x"4120", x"4177",
        x"41CD", x"4223", x"4279", x"42CF", x"4325", x"437A", x"43D0", x"4425",
        x"447A", x"44CF", x"4523", x"4578", x"45CC", x"4620", x"4674", x"46C8",
        x"471C", x"476F", x"47C3", x"4816", x"4869", x"48BC", x"490E", x"4961",
        x"49B3", x"4A05", x"4A57", x"4AA9", x"4AFA", x"4B4C", x"4B9D", x"4BEE",
        x"4C3F", x"4C8F", x"4CE0", x"4D30", x"4D80", x"4DD0", x"4E20", x"4E6F",
        x"4EBF", x"4F0E", x"4F5D", x"4FAC", x"4FFA", x"5049", x"5097", x"50E5",
        x"5133", x"5180", x"51CE", x"521B", x"5268", x"52B5", x"5301", x"534E",
        x"539A", x"53E6", x"5432", x"547D", x"54C9", x"5514", x"555F", x"55AA",
        x"55F4", x"563F", x"5689", x"56D3", x"571D", x"5766", x"57B0", x"57F9",
        x"5842", x"588A", x"58D3", x"591B", x"5963", x"59AB", x"59F3", x"5A3A",
        x"5A81", x"5AC8", x"5B0F", x"5B56", x"5B9C", x"5BE2", x"5C28", x"5C6D",
        x"5CB3", x"5CF8", x"5D3D", x"5D82", x"5DC6", x"5E0B", x"5E4F", x"5E93",
        x"5ED6", x"5F1A", x"5F5D", x"5FA0", x"5FE2", x"6025", x"6067", x"60A9",
        x"60EB", x"612D", x"616E", x"61AF", x"61F0", x"6230", x"6271", x"62B1",
        x"62F1", x"6330", x"6370", x"63AF", x"63EE", x"642D", x"646B", x"64A9",
        x"64E7", x"6525", x"6562", x"65A0", x"65DD", x"6619", x"6656", x"6692",
        x"66CE", x"670A", x"6745", x"6781", x"67BC", x"67F7", x"6831", x"686B",
        x"68A5", x"68DF", x"6919", x"6952", x"698B", x"69C4", x"69FC", x"6A34",
        x"6A6C", x"6AA4", x"6ADB", x"6B13", x"6B4A", x"6B80", x"6BB7", x"6BED",
        x"6C23", x"6C58", x"6C8E", x"6CC3", x"6CF8", x"6D2C", x"6D61", x"6D95",
        x"6DC9", x"6DFC", x"6E30", x"6E63", x"6E95", x"6EC8", x"6EFA", x"6F2C",
        x"6F5E", x"6F8F", x"6FC0", x"6FF1", x"7022", x"7052", x"7082", x"70B2",
        x"70E1", x"7111", x"7140", x"716E", x"719D", x"71CB", x"71F9", x"7226",
        x"7254", x"7281", x"72AE", x"72DA", x"7306", x"7332", x"735E", x"7389",
        x"73B5", x"73DF", x"740A", x"7434", x"745E", x"7488", x"74B1", x"74DB",
        x"7503", x"752C", x"7554", x"757C", x"75A4", x"75CC", x"75F3", x"761A",
        x"7640", x"7667", x"768D", x"76B2", x"76D8", x"76FD", x"7722", x"7747",
        x"776B", x"778F", x"77B3", x"77D6", x"77F9", x"781C", x"783F", x"7861",
        x"7883", x"78A5", x"78C6", x"78E7", x"7908", x"7929", x"7949", x"7969",
        x"7989", x"79A8", x"79C7", x"79E6", x"7A04", x"7A23", x"7A41", x"7A5E",
        x"7A7C", x"7A99", x"7AB5", x"7AD2", x"7AEE", x"7B0A", x"7B25", x"7B41",
        x"7B5C", x"7B76", x"7B91", x"7BAB", x"7BC4", x"7BDE", x"7BF7", x"7C10",
        x"7C29", x"7C41", x"7C59", x"7C70", x"7C88", x"7C9F", x"7CB6", x"7CCC",
        x"7CE2", x"7CF8", x"7D0E", x"7D23", x"7D38", x"7D4D", x"7D61", x"7D75",
        x"7D89", x"7D9C", x"7DB0", x"7DC2", x"7DD5", x"7DE7", x"7DF9", x"7E0B",
        x"7E1C", x"7E2D", x"7E3E", x"7E4E", x"7E5E", x"7E6E", x"7E7E", x"7E8D",
        x"7E9C", x"7EAA", x"7EB9", x"7EC7", x"7ED4", x"7EE2", x"7EEF", x"7EFC",
        x"7F08", x"7F14", x"7F20", x"7F2C", x"7F37", x"7F42", x"7F4C", x"7F57",
        x"7F61", x"7F6A", x"7F74", x"7F7D", x"7F86", x"7F8E", x"7F96", x"7F9E",
        x"7FA6", x"7FAD", x"7FB4", x"7FBB", x"7FC1", x"7FC7", x"7FCD", x"7FD2",
        x"7FD7", x"7FDC", x"7FE0", x"7FE4", x"7FE8", x"7FEC", x"7FEF", x"7FF2",
        x"7FF5", x"7FF7", x"7FF9", x"7FFB", x"7FFC", x"7FFD", x"7FFE", x"7FFE",
        x"7FFF", x"7FFE", x"7FFE", x"7FFD", x"7FFC", x"7FFB", x"7FF9", x"7FF7",
        x"7FF5", x"7FF2", x"7FEF", x"7FEC", x"7FE8", x"7FE4", x"7FE0", x"7FDC",
        x"7FD7", x"7FD2", x"7FCD", x"7FC7", x"7FC1", x"7FBB", x"7FB4", x"7FAD",
        x"7FA6", x"7F9E", x"7F96", x"7F8E", x"7F86", x"7F7D", x"7F74", x"7F6A",
        x"7F61", x"7F57", x"7F4C", x"7F42", x"7F37", x"7F2C", x"7F20", x"7F14",
        x"7F08", x"7EFC", x"7EEF", x"7EE2", x"7ED4", x"7EC7", x"7EB9", x"7EAA",
        x"7E9C", x"7E8D", x"7E7E", x"7E6E", x"7E5E", x"7E4E", x"7E3E", x"7E2D",
        x"7E1C", x"7E0B", x"7DF9", x"7DE7", x"7DD5", x"7DC2", x"7DB0", x"7D9C",
        x"7D89", x"7D75", x"7D61", x"7D4D", x"7D38", x"7D23", x"7D0E", x"7CF8",
        x"7CE2", x"7CCC", x"7CB6", x"7C9F", x"7C88", x"7C70", x"7C59", x"7C41",
        x"7C29", x"7C10", x"7BF7", x"7BDE", x"7BC4", x"7BAB", x"7B91", x"7B76",
        x"7B5C", x"7B41", x"7B25", x"7B0A", x"7AEE", x"7AD2", x"7AB5", x"7A99",
        x"7A7C", x"7A5E", x"7A41", x"7A23", x"7A04", x"79E6", x"79C7", x"79A8",
        x"7989", x"7969", x"7949", x"7929", x"7908", x"78E7", x"78C6", x"78A5",
        x"7883", x"7861", x"783F", x"781C", x"77F9", x"77D6", x"77B3", x"778F",
        x"776B", x"7747", x"7722", x"76FD", x"76D8", x"76B2", x"768D", x"7667",
        x"7640", x"761A", x"75F3", x"75CC", x"75A4", x"757C", x"7554", x"752C",
        x"7503", x"74DB", x"74B1", x"7488", x"745E", x"7434", x"740A", x"73DF",
        x"73B5", x"7389", x"735E", x"7332", x"7306", x"72DA", x"72AE", x"7281",
        x"7254", x"7226", x"71F9", x"71CB", x"719D", x"716E", x"7140", x"7111",
        x"70E1", x"70B2", x"7082", x"7052", x"7022", x"6FF1", x"6FC0", x"6F8F",
        x"6F5E", x"6F2C", x"6EFA", x"6EC8", x"6E95", x"6E63", x"6E30", x"6DFC",
        x"6DC9", x"6D95", x"6D61", x"6D2C", x"6CF8", x"6CC3", x"6C8E", x"6C58",
        x"6C23", x"6BED", x"6BB7", x"6B80", x"6B4A", x"6B13", x"6ADB", x"6AA4",
        x"6A6C", x"6A34", x"69FC", x"69C4", x"698B", x"6952", x"6919", x"68DF",
        x"68A5", x"686B", x"6831", x"67F7", x"67BC", x"6781", x"6745", x"670A",
        x"66CE", x"6692", x"6656", x"6619", x"65DD", x"65A0", x"6562", x"6525",
        x"64E7", x"64A9", x"646B", x"642D", x"63EE", x"63AF", x"6370", x"6330",
        x"62F1", x"62B1", x"6271", x"6230", x"61F0", x"61AF", x"616E", x"612D",
        x"60EB", x"60A9", x"6067", x"6025", x"5FE2", x"5FA0", x"5F5D", x"5F1A",
        x"5ED6", x"5E93", x"5E4F", x"5E0B", x"5DC6", x"5D82", x"5D3D", x"5CF8",
        x"5CB3", x"5C6D", x"5C28", x"5BE2", x"5B9C", x"5B56", x"5B0F", x"5AC8",
        x"5A81", x"5A3A", x"59F3", x"59AB", x"5963", x"591B", x"58D3", x"588A",
        x"5842", x"57F9", x"57B0", x"5766", x"571D", x"56D3", x"5689", x"563F",
        x"55F4", x"55AA", x"555F", x"5514", x"54C9", x"547D", x"5432", x"53E6",
        x"539A", x"534E", x"5301", x"52B5", x"5268", x"521B", x"51CE", x"5180",
        x"5133", x"50E5", x"5097", x"5049", x"4FFA", x"4FAC", x"4F5D", x"4F0E",
        x"4EBF", x"4E6F", x"4E20", x"4DD0", x"4D80", x"4D30", x"4CE0", x"4C8F",
        x"4C3F", x"4BEE", x"4B9D", x"4B4C", x"4AFA", x"4AA9", x"4A57", x"4A05",
        x"49B3", x"4961", x"490E", x"48BC", x"4869", x"4816", x"47C3", x"476F",
        x"471C", x"46C8", x"4674", x"4620", x"45CC", x"4578", x"4523", x"44CF",
        x"447A", x"4425", x"43D0", x"437A", x"4325", x"42CF", x"4279", x"4223",
        x"41CD", x"4177", x"4120", x"40CA", x"4073", x"401C", x"3FC5", x"3F6E",
        x"3F16", x"3EBF", x"3E67", x"3E0F", x"3DB7", x"3D5F", x"3D07", x"3CAE",
        x"3C56", x"3BFD", x"3BA4", x"3B4B", x"3AF2", x"3A99", x"3A3F", x"39E6",
        x"398C", x"3932", x"38D8", x"387E", x"3824", x"37C9", x"376F", x"3714",
        x"36B9", x"365E", x"3603", x"35A8", x"354D", x"34F1", x"3496", x"343A",
        x"33DE", x"3382", x"3326", x"32CA", x"326D", x"3211", x"31B4", x"3158",
        x"30FB", x"309E", x"3041", x"2FE4", x"2F86", x"2F29", x"2ECC", x"2E6E",
        x"2E10", x"2DB2", x"2D54", x"2CF6", x"2C98", x"2C3A", x"2BDB", x"2B7D",
        x"2B1E", x"2AC0", x"2A61", x"2A02", x"29A3", x"2944", x"28E5", x"2885",
        x"2826", x"27C6", x"2767", x"2707", x"26A7", x"2647", x"25E7", x"2587",
        x"2527", x"24C7", x"2467", x"2406", x"23A6", x"2345", x"22E4", x"2284",
        x"2223", x"21C2", x"2161", x"2100", x"209F", x"203D", x"1FDC", x"1F7B",
        x"1F19", x"1EB8", x"1E56", x"1DF4", x"1D93", x"1D31", x"1CCF", x"1C6D",
        x"1C0B", x"1BA9", x"1B46", x"1AE4", x"1A82", x"1A20", x"19BD", x"195B",
        x"18F8", x"1895", x"1833", x"17D0", x"176D", x"170A", x"16A7", x"1644",
        x"15E1", x"157E", x"151B", x"14B8", x"1455", x"13F2", x"138E", x"132B",
        x"12C7", x"1264", x"1200", x"119D", x"1139", x"10D6", x"1072", x"100E",
        x"0FAB", x"0F47", x"0EE3", x"0E7F", x"0E1B", x"0DB7", x"0D53", x"0CEF",
        x"0C8B", x"0C27", x"0BC3", x"0B5F", x"0AFB", x"0A97", x"0A32", x"09CE",
        x"096A", x"0906", x"08A1", x"083D", x"07D9", x"0774", x"0710", x"06AC",
        x"0647", x"05E3", x"057E", x"051A", x"04B6", x"0451", x"03ED", x"0388",
        x"0324", x"02BF", x"025B", x"01F6", x"0192", x"012D", x"00C9", x"0064",
        x"0000", x"FF9C", x"FF37", x"FED3", x"FE6E", x"FE0A", x"FDA5", x"FD41",
        x"FCDC", x"FC78", x"FC13", x"FBAF", x"FB4A", x"FAE6", x"FA82", x"FA1D",
        x"F9B9", x"F954", x"F8F0", x"F88C", x"F827", x"F7C3", x"F75F", x"F6FA",
        x"F696", x"F632", x"F5CE", x"F569", x"F505", x"F4A1", x"F43D", x"F3D9",
        x"F375", x"F311", x"F2AD", x"F249", x"F1E5", x"F181", x"F11D", x"F0B9",
        x"F055", x"EFF2", x"EF8E", x"EF2A", x"EEC7", x"EE63", x"EE00", x"ED9C",
        x"ED39", x"ECD5", x"EC72", x"EC0E", x"EBAB", x"EB48", x"EAE5", x"EA82",
        x"EA1F", x"E9BC", x"E959", x"E8F6", x"E893", x"E830", x"E7CD", x"E76B",
        x"E708", x"E6A5", x"E643", x"E5E0", x"E57E", x"E51C", x"E4BA", x"E457",
        x"E3F5", x"E393", x"E331", x"E2CF", x"E26D", x"E20C", x"E1AA", x"E148",
        x"E0E7", x"E085", x"E024", x"DFC3", x"DF61", x"DF00", x"DE9F", x"DE3E",
        x"DDDD", x"DD7C", x"DD1C", x"DCBB", x"DC5A", x"DBFA", x"DB99", x"DB39",
        x"DAD9", x"DA79", x"DA19", x"D9B9", x"D959", x"D8F9", x"D899", x"D83A",
        x"D7DA", x"D77B", x"D71B", x"D6BC", x"D65D", x"D5FE", x"D59F", x"D540",
        x"D4E2", x"D483", x"D425", x"D3C6", x"D368", x"D30A", x"D2AC", x"D24E",
        x"D1F0", x"D192", x"D134", x"D0D7", x"D07A", x"D01C", x"CFBF", x"CF62",
        x"CF05", x"CEA8", x"CE4C", x"CDEF", x"CD93", x"CD36", x"CCDA", x"CC7E",
        x"CC22", x"CBC6", x"CB6A", x"CB0F", x"CAB3", x"CA58", x"C9FD", x"C9A2",
        x"C947", x"C8EC", x"C891", x"C837", x"C7DC", x"C782", x"C728", x"C6CE",
        x"C674", x"C61A", x"C5C1", x"C567", x"C50E", x"C4B5", x"C45C", x"C403",
        x"C3AA", x"C352", x"C2F9", x"C2A1", x"C249", x"C1F1", x"C199", x"C141",
        x"C0EA", x"C092", x"C03B", x"BFE4", x"BF8D", x"BF36", x"BEE0", x"BE89",
        x"BE33", x"BDDD", x"BD87", x"BD31", x"BCDB", x"BC86", x"BC30", x"BBDB",
        x"BB86", x"BB31", x"BADD", x"BA88", x"BA34", x"B9E0", x"B98C", x"B938",
        x"B8E4", x"B891", x"B83D", x"B7EA", x"B797", x"B744", x"B6F2", x"B69F",
        x"B64D", x"B5FB", x"B5A9", x"B557", x"B506", x"B4B4", x"B463", x"B412",
        x"B3C1", x"B371", x"B320", x"B2D0", x"B280", x"B230", x"B1E0", x"B191",
        x"B141", x"B0F2", x"B0A3", x"B054", x"B006", x"AFB7", x"AF69", x"AF1B",
        x"AECD", x"AE80", x"AE32", x"ADE5", x"AD98", x"AD4B", x"ACFF", x"ACB2",
        x"AC66", x"AC1A", x"ABCE", x"AB83", x"AB37", x"AAEC", x"AAA1", x"AA56",
        x"AA0C", x"A9C1", x"A977", x"A92D", x"A8E3", x"A89A", x"A850", x"A807",
        x"A7BE", x"A776", x"A72D", x"A6E5", x"A69D", x"A655", x"A60D", x"A5C6",
        x"A57F", x"A538", x"A4F1", x"A4AA", x"A464", x"A41E", x"A3D8", x"A393",
        x"A34D", x"A308", x"A2C3", x"A27E", x"A23A", x"A1F5", x"A1B1", x"A16D",
        x"A12A", x"A0E6", x"A0A3", x"A060", x"A01E", x"9FDB", x"9F99", x"9F57",
        x"9F15", x"9ED3", x"9E92", x"9E51", x"9E10", x"9DD0", x"9D8F", x"9D4F",
        x"9D0F", x"9CD0", x"9C90", x"9C51", x"9C12", x"9BD3", x"9B95", x"9B57",
        x"9B19", x"9ADB", x"9A9E", x"9A60", x"9A23", x"99E7", x"99AA", x"996E",
        x"9932", x"98F6", x"98BB", x"987F", x"9844", x"9809", x"97CF", x"9795",
        x"975B", x"9721", x"96E7", x"96AE", x"9675", x"963C", x"9604", x"95CC",
        x"9594", x"955C", x"9525", x"94ED", x"94B6", x"9480", x"9449", x"9413",
        x"93DD", x"93A8", x"9372", x"933D", x"9308", x"92D4", x"929F", x"926B",
        x"9237", x"9204", x"91D0", x"919D", x"916B", x"9138", x"9106", x"90D4",
        x"90A2", x"9071", x"9040", x"900F", x"8FDE", x"8FAE", x"8F7E", x"8F4E",
        x"8F1F", x"8EEF", x"8EC0", x"8E92", x"8E63", x"8E35", x"8E07", x"8DDA",
        x"8DAC", x"8D7F", x"8D52", x"8D26", x"8CFA", x"8CCE", x"8CA2", x"8C77",
        x"8C4B", x"8C21", x"8BF6", x"8BCC", x"8BA2", x"8B78", x"8B4F", x"8B25",
        x"8AFD", x"8AD4", x"8AAC", x"8A84", x"8A5C", x"8A34", x"8A0D", x"89E6",
        x"89C0", x"8999", x"8973", x"894E", x"8928", x"8903", x"88DE", x"88B9",
        x"8895", x"8871", x"884D", x"882A", x"8807", x"87E4", x"87C1", x"879F",
        x"877D", x"875B", x"873A", x"8719", x"86F8", x"86D7", x"86B7", x"8697",
        x"8677", x"8658", x"8639", x"861A", x"85FC", x"85DD", x"85BF", x"85A2",
        x"8584", x"8567", x"854B", x"852E", x"8512", x"84F6", x"84DB", x"84BF",
        x"84A4", x"848A", x"846F", x"8455", x"843C", x"8422", x"8409", x"83F0",
        x"83D7", x"83BF", x"83A7", x"8390", x"8378", x"8361", x"834A", x"8334",
        x"831E", x"8308", x"82F2", x"82DD", x"82C8", x"82B3", x"829F", x"828B",
        x"8277", x"8264", x"8250", x"823E", x"822B", x"8219", x"8207", x"81F5",
        x"81E4", x"81D3", x"81C2", x"81B2", x"81A2", x"8192", x"8182", x"8173",
        x"8164", x"8156", x"8147", x"8139", x"812C", x"811E", x"8111", x"8104",
        x"80F8", x"80EC", x"80E0", x"80D4", x"80C9", x"80BE", x"80B4", x"80A9",
        x"809F", x"8096", x"808C", x"8083", x"807A", x"8072", x"806A", x"8062",
        x"805A", x"8053", x"804C", x"8045", x"803F", x"8039", x"8033", x"802E",
        x"8029", x"8024", x"8020", x"801C", x"8018", x"8014", x"8011", x"800E",
        x"800B", x"8009", x"8007", x"8005", x"8004", x"8003", x"8002", x"8002",
        x"8001", x"8002", x"8002", x"8003", x"8004", x"8005", x"8007", x"8009",
        x"800B", x"800E", x"8011", x"8014", x"8018", x"801C", x"8020", x"8024",
        x"8029", x"802E", x"8033", x"8039", x"803F", x"8045", x"804C", x"8053",
        x"805A", x"8062", x"806A", x"8072", x"807A", x"8083", x"808C", x"8096",
        x"809F", x"80A9", x"80B4", x"80BE", x"80C9", x"80D4", x"80E0", x"80EC",
        x"80F8", x"8104", x"8111", x"811E", x"812C", x"8139", x"8147", x"8156",
        x"8164", x"8173", x"8182", x"8192", x"81A2", x"81B2", x"81C2", x"81D3",
        x"81E4", x"81F5", x"8207", x"8219", x"822B", x"823E", x"8250", x"8264",
        x"8277", x"828B", x"829F", x"82B3", x"82C8", x"82DD", x"82F2", x"8308",
        x"831E", x"8334", x"834A", x"8361", x"8378", x"8390", x"83A7", x"83BF",
        x"83D7", x"83F0", x"8409", x"8422", x"843C", x"8455", x"846F", x"848A",
        x"84A4", x"84BF", x"84DB", x"84F6", x"8512", x"852E", x"854B", x"8567",
        x"8584", x"85A2", x"85BF", x"85DD", x"85FC", x"861A", x"8639", x"8658",
        x"8677", x"8697", x"86B7", x"86D7", x"86F8", x"8719", x"873A", x"875B",
        x"877D", x"879F", x"87C1", x"87E4", x"8807", x"882A", x"884D", x"8871",
        x"8895", x"88B9", x"88DE", x"8903", x"8928", x"894E", x"8973", x"8999",
        x"89C0", x"89E6", x"8A0D", x"8A34", x"8A5C", x"8A84", x"8AAC", x"8AD4",
        x"8AFD", x"8B25", x"8B4F", x"8B78", x"8BA2", x"8BCC", x"8BF6", x"8C21",
        x"8C4B", x"8C77", x"8CA2", x"8CCE", x"8CFA", x"8D26", x"8D52", x"8D7F",
        x"8DAC", x"8DDA", x"8E07", x"8E35", x"8E63", x"8E92", x"8EC0", x"8EEF",
        x"8F1F", x"8F4E", x"8F7E", x"8FAE", x"8FDE", x"900F", x"9040", x"9071",
        x"90A2", x"90D4", x"9106", x"9138", x"916B", x"919D", x"91D0", x"9204",
        x"9237", x"926B", x"929F", x"92D4", x"9308", x"933D", x"9372", x"93A8",
        x"93DD", x"9413", x"9449", x"9480", x"94B6", x"94ED", x"9525", x"955C",
        x"9594", x"95CC", x"9604", x"963C", x"9675", x"96AE", x"96E7", x"9721",
        x"975B", x"9795", x"97CF", x"9809", x"9844", x"987F", x"98BB", x"98F6",
        x"9932", x"996E", x"99AA", x"99E7", x"9A23", x"9A60", x"9A9E", x"9ADB",
        x"9B19", x"9B57", x"9B95", x"9BD3", x"9C12", x"9C51", x"9C90", x"9CD0",
        x"9D0F", x"9D4F", x"9D8F", x"9DD0", x"9E10", x"9E51", x"9E92", x"9ED3",
        x"9F15", x"9F57", x"9F99", x"9FDB", x"A01E", x"A060", x"A0A3", x"A0E6",
        x"A12A", x"A16D", x"A1B1", x"A1F5", x"A23A", x"A27E", x"A2C3", x"A308",
        x"A34D", x"A393", x"A3D8", x"A41E", x"A464", x"A4AA", x"A4F1", x"A538",
        x"A57F", x"A5C6", x"A60D", x"A655", x"A69D", x"A6E5", x"A72D", x"A776",
        x"A7BE", x"A807", x"A850", x"A89A", x"A8E3", x"A92D", x"A977", x"A9C1",
        x"AA0C", x"AA56", x"AAA1", x"AAEC", x"AB37", x"AB83", x"ABCE", x"AC1A",
        x"AC66", x"ACB2", x"ACFF", x"AD4B", x"AD98", x"ADE5", x"AE32", x"AE80",
        x"AECD", x"AF1B", x"AF69", x"AFB7", x"B006", x"B054", x"B0A3", x"B0F2",
        x"B141", x"B191", x"B1E0", x"B230", x"B280", x"B2D0", x"B320", x"B371",
        x"B3C1", x"B412", x"B463", x"B4B4", x"B506", x"B557", x"B5A9", x"B5FB",
        x"B64D", x"B69F", x"B6F2", x"B744", x"B797", x"B7EA", x"B83D", x"B891",
        x"B8E4", x"B938", x"B98C", x"B9E0", x"BA34", x"BA88", x"BADD", x"BB31",
        x"BB86", x"BBDB", x"BC30", x"BC86", x"BCDB", x"BD31", x"BD87", x"BDDD",
        x"BE33", x"BE89", x"BEE0", x"BF36", x"BF8D", x"BFE4", x"C03B", x"C092",
        x"C0EA", x"C141", x"C199", x"C1F1", x"C249", x"C2A1", x"C2F9", x"C352",
        x"C3AA", x"C403", x"C45C", x"C4B5", x"C50E", x"C567", x"C5C1", x"C61A",
        x"C674", x"C6CE", x"C728", x"C782", x"C7DC", x"C837", x"C891", x"C8EC",
        x"C947", x"C9A2", x"C9FD", x"CA58", x"CAB3", x"CB0F", x"CB6A", x"CBC6",
        x"CC22", x"CC7E", x"CCDA", x"CD36", x"CD93", x"CDEF", x"CE4C", x"CEA8",
        x"CF05", x"CF62", x"CFBF", x"D01C", x"D07A", x"D0D7", x"D134", x"D192",
        x"D1F0", x"D24E", x"D2AC", x"D30A", x"D368", x"D3C6", x"D425", x"D483",
        x"D4E2", x"D540", x"D59F", x"D5FE", x"D65D", x"D6BC", x"D71B", x"D77B",
        x"D7DA", x"D83A", x"D899", x"D8F9", x"D959", x"D9B9", x"DA19", x"DA79",
        x"DAD9", x"DB39", x"DB99", x"DBFA", x"DC5A", x"DCBB", x"DD1C", x"DD7C",
        x"DDDD", x"DE3E", x"DE9F", x"DF00", x"DF61", x"DFC3", x"E024", x"E085",
        x"E0E7", x"E148", x"E1AA", x"E20C", x"E26D", x"E2CF", x"E331", x"E393",
        x"E3F5", x"E457", x"E4BA", x"E51C", x"E57E", x"E5E0", x"E643", x"E6A5",
        x"E708", x"E76B", x"E7CD", x"E830", x"E893", x"E8F6", x"E959", x"E9BC",
        x"EA1F", x"EA82", x"EAE5", x"EB48", x"EBAB", x"EC0E", x"EC72", x"ECD5",
        x"ED39", x"ED9C", x"EE00", x"EE63", x"EEC7", x"EF2A", x"EF8E", x"EFF2",
        x"F055", x"F0B9", x"F11D", x"F181", x"F1E5", x"F249", x"F2AD", x"F311",
        x"F375", x"F3D9", x"F43D", x"F4A1", x"F505", x"F569", x"F5CE", x"F632",
        x"F696", x"F6FA", x"F75F", x"F7C3", x"F827", x"F88C", x"F8F0", x"F954",
        x"F9B9", x"FA1D", x"FA82", x"FAE6", x"FB4A", x"FBAF", x"FC13", x"FC78",
        x"FCDC", x"FD41", x"FDA5", x"FE0A", x"FE6E", x"FED3", x"FF37", x"FF9C"
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            dout <= lut(to_integer(unsigned(addr)));
        end if;
    end process;
end arch;