Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity guitar_lut is
    generic (
        DEPTH : integer := 2048;
        WIDTH : integer := 16
    );
    port (
        clk   : in  std_logic;
        addr  : in  std_logic_vector(10 downto 0);
        dout  : out std_logic_vector(WIDTH-1 downto 0)
    );
end guitar_lut;

architecture arch of guitar_lut is
    type lut_array is array(0 to DEPTH-1) of std_logic_vector(WIDTH-1 downto 0);
    signal lut: lut_array := (
x"0000",
x"028C",
x"0519",
x"07A5",
x"0A31",
x"0CBC",
x"0F46",
x"11CF",
x"1458",
x"16DE",
x"1964",
x"1BE7",
x"1E69",
x"20E9",
x"2367",
x"25E3",
x"285C",
x"2AD2",
x"2D46",
x"2FB7",
x"3225",
x"3490",
x"36F7",
x"395B",
x"3BBC",
x"3E18",
x"4071",
x"42C5",
x"4516",
x"4762",
x"49AA",
x"4BED",
x"4E2B",
x"5065",
x"529A",
x"54C9",
x"56F4",
x"5919",
x"5B39",
x"5D53",
x"5F68",
x"6177",
x"6380",
x"6584",
x"6781",
x"6978",
x"6B69",
x"6D54",
x"6F38",
x"7116",
x"72EE",
x"74BF",
x"7689",
x"784D",
x"7A0A",
x"7BC0",
x"7D6F",
x"7F17",
x"80B9",
x"8253",
x"83E6",
x"8572",
x"86F8",
x"8875",
x"89EC",
x"8B5C",
x"8CC4",
x"8E25",
x"8F7E",
x"90D1",
x"921C",
x"9360",
x"949C",
x"95D1",
x"96FF",
x"9826",
x"9945",
x"9A5D",
x"9B6E",
x"9C78",
x"9D7A",
x"9E76",
x"9F6A",
x"A057",
x"A13D",
x"A21B",
x"A2F3",
x"A3C4",
x"A48E",
x"A551",
x"A60E",
x"A6C3",
x"A772",
x"A81A",
x"A8BC",
x"A957",
x"A9EB",
x"AA79",
x"AB01",
x"AB83",
x"ABFE",
x"AC74",
x"ACE3",
x"AD4C",
x"ADB0",
x"AE0D",
x"AE65",
x"AEB7",
x"AF04",
x"AF4C",
x"AF8E",
x"AFCA",
x"B002",
x"B034",
x"B062",
x"B08A",
x"B0AE",
x"B0CD",
x"B0E7",
x"B0FD",
x"B10F",
x"B11C",
x"B125",
x"B12A",
x"B12A",
x"B127",
x"B120",
x"B116",
x"B108",
x"B0F6",
x"B0E1",
x"B0C8",
x"B0AD",
x"B08E",
x"B06C",
x"B047",
x"B020",
x"AFF6",
x"AFC9",
x"AF99",
x"AF68",
x"AF33",
x"AEFD",
x"AEC5",
x"AE8A",
x"AE4E",
x"AE0F",
x"ADCF",
x"AD8D",
x"AD4A",
x"AD05",
x"ACBF",
x"AC77",
x"AC2E",
x"ABE4",
x"AB99",
x"AB4D",
x"AB00",
x"AAB2",
x"AA63",
x"AA13",
x"A9C3",
x"A973",
x"A922",
x"A8D0",
x"A87E",
x"A82C",
x"A7DA",
x"A787",
x"A734",
x"A6E1",
x"A68F",
x"A63C",
x"A5E9",
x"A597",
x"A544",
x"A4F2",
x"A4A1",
x"A44F",
x"A3FE",
x"A3AE",
x"A35D",
x"A30E",
x"A2BF",
x"A270",
x"A222",
x"A1D5",
x"A188",
x"A13C",
x"A0F1",
x"A0A6",
x"A05C",
x"A013",
x"9FCB",
x"9F83",
x"9F3C",
x"9EF7",
x"9EB1",
x"9E6D",
x"9E2A",
x"9DE7",
x"9DA6",
x"9D65",
x"9D25",
x"9CE6",
x"9CA8",
x"9C6B",
x"9C2F",
x"9BF3",
x"9BB9",
x"9B7F",
x"9B46",
x"9B0E",
x"9AD7",
x"9AA1",
x"9A6B",
x"9A36",
x"9A02",
x"99CF",
x"999D",
x"996C",
x"993B",
x"990B",
x"98DB",
x"98AD",
x"987F",
x"9851",
x"9825",
x"97F9",
x"97CD",
x"97A2",
x"9778",
x"974E",
x"9725",
x"96FC",
x"96D4",
x"96AC",
x"9685",
x"965E",
x"9638",
x"9611",
x"95EB",
x"95C6",
x"95A1",
x"957C",
x"9557",
x"9533",
x"950E",
x"94EA",
x"94C7",
x"94A3",
x"947F",
x"945C",
x"9438",
x"9415",
x"93F2",
x"93CE",
x"93AB",
x"9388",
x"9365",
x"9341",
x"931E",
x"92FA",
x"92D7",
x"92B3",
x"928F",
x"926B",
x"9247",
x"9223",
x"91FE",
x"91DA",
x"91B5",
x"9190",
x"916A",
x"9145",
x"911F",
x"90F9",
x"90D3",
x"90AC",
x"9085",
x"905E",
x"9036",
x"900E",
x"8FE6",
x"8FBE",
x"8F95",
x"8F6C",
x"8F42",
x"8F19",
x"8EEF",
x"8EC4",
x"8E99",
x"8E6E",
x"8E43",
x"8E17",
x"8DEB",
x"8DBF",
x"8D92",
x"8D65",
x"8D38",
x"8D0A",
x"8CDC",
x"8CAE",
x"8C80",
x"8C51",
x"8C22",
x"8BF2",
x"8BC3",
x"8B93",
x"8B62",
x"8B32",
x"8B01",
x"8AD0",
x"8A9F",
x"8A6E",
x"8A3D",
x"8A0B",
x"89D9",
x"89A7",
x"8975",
x"8942",
x"8910",
x"88DD",
x"88AA",
x"8877",
x"8844",
x"8811",
x"87DE",
x"87AA",
x"8777",
x"8744",
x"8710",
x"86DD",
x"86A9",
x"8676",
x"8642",
x"860F",
x"85DB",
x"85A8",
x"8574",
x"8541",
x"850E",
x"84DA",
x"84A7",
x"8474",
x"8441",
x"840E",
x"83DB",
x"83A8",
x"8376",
x"8343",
x"8311",
x"82DF",
x"82AD",
x"827B",
x"8249",
x"8217",
x"81E6",
x"81B5",
x"8184",
x"8153",
x"8122",
x"80F1",
x"80C1",
x"8091",
x"8061",
x"8031",
x"8001",
x"7FD2",
x"7FA2",
x"7F73",
x"7F45",
x"7F16",
x"7EE7",
x"7EB9",
x"7E8B",
x"7E5D",
x"7E2F",
x"7E02",
x"7DD4",
x"7DA7",
x"7D7A",
x"7D4D",
x"7D20",
x"7CF4",
x"7CC7",
x"7C9B",
x"7C6F",
x"7C43",
x"7C17",
x"7BEB",
x"7BC0",
x"7B94",
x"7B69",
x"7B3E",
x"7B13",
x"7AE7",
x"7ABC",
x"7A91",
x"7A67",
x"7A3C",
x"7A11",
x"79E6",
x"79BC",
x"7991",
x"7966",
x"793C",
x"7911",
x"78E7",
x"78BC",
x"7891",
x"7867",
x"783C",
x"7811",
x"77E6",
x"77BC",
x"7791",
x"7766",
x"773B",
x"7710",
x"76E4",
x"76B9",
x"768E",
x"7662",
x"7636",
x"760B",
x"75DF",
x"75B3",
x"7587",
x"755A",
x"752E",
x"7501",
x"74D4",
x"74A7",
x"747A",
x"744D",
x"741F",
x"73F2",
x"73C4",
x"7396",
x"7368",
x"7339",
x"730B",
x"72DC",
x"72AD",
x"727D",
x"724E",
x"721E",
x"71EF",
x"71BF",
x"718E",
x"715E",
x"712D",
x"70FC",
x"70CB",
x"709A",
x"7069",
x"7037",
x"7005",
x"6FD3",
x"6FA1",
x"6F6F",
x"6F3C",
x"6F0A",
x"6ED7",
x"6EA4",
x"6E71",
x"6E3D",
x"6E0A",
x"6DD6",
x"6DA3",
x"6D6F",
x"6D3B",
x"6D07",
x"6CD3",
x"6C9E",
x"6C6A",
x"6C35",
x"6C01",
x"6BCC",
x"6B97",
x"6B63",
x"6B2E",
x"6AF9",
x"6AC4",
x"6A8F",
x"6A5A",
x"6A26",
x"69F1",
x"69BC",
x"6987",
x"6952",
x"691D",
x"68E8",
x"68B4",
x"687F",
x"684B",
x"6816",
x"67E2",
x"67AD",
x"6779",
x"6745",
x"6711",
x"66DD",
x"66A9",
x"6676",
x"6642",
x"660F",
x"65DC",
x"65A9",
x"6577",
x"6544",
x"6512",
x"64E0",
x"64AE",
x"647C",
x"644A",
x"6419",
x"63E8",
x"63B7",
x"6387",
x"6356",
x"6326",
x"62F7",
x"62C7",
x"6298",
x"6269",
x"623A",
x"620B",
x"61DD",
x"61AF",
x"6182",
x"6154",
x"6127",
x"60FA",
x"60CE",
x"60A2",
x"6076",
x"604A",
x"601E",
x"5FF3",
x"5FC8",
x"5F9E",
x"5F73",
x"5F49",
x"5F20",
x"5EF6",
x"5ECD",
x"5EA4",
x"5E7B",
x"5E53",
x"5E2A",
x"5E02",
x"5DDA",
x"5DB3",
x"5D8C",
x"5D64",
x"5D3E",
x"5D17",
x"5CF0",
x"5CCA",
x"5CA4",
x"5C7E",
x"5C58",
x"5C32",
x"5C0D",
x"5BE8",
x"5BC2",
x"5B9D",
x"5B78",
x"5B54",
x"5B2F",
x"5B0A",
x"5AE6",
x"5AC1",
x"5A9D",
x"5A78",
x"5A54",
x"5A30",
x"5A0B",
x"59E7",
x"59C3",
x"599F",
x"597A",
x"5956",
x"5932",
x"590D",
x"58E9",
x"58C4",
x"58A0",
x"587B",
x"5856",
x"5831",
x"580C",
x"57E7",
x"57C2",
x"579C",
x"5777",
x"5751",
x"572B",
x"5705",
x"56DF",
x"56B8",
x"5691",
x"566A",
x"5643",
x"561C",
x"55F4",
x"55CC",
x"55A4",
x"557C",
x"5553",
x"552A",
x"5501",
x"54D7",
x"54AE",
x"5484",
x"5459",
x"542E",
x"5403",
x"53D8",
x"53AC",
x"5380",
x"5354",
x"5328",
x"52FB",
x"52CD",
x"52A0",
x"5272",
x"5243",
x"5215",
x"51E6",
x"51B6",
x"5187",
x"5156",
x"5126",
x"50F5",
x"50C4",
x"5093",
x"5061",
x"502F",
x"4FFC",
x"4FCA",
x"4F97",
x"4F63",
x"4F2F",
x"4EFB",
x"4EC7",
x"4E92",
x"4E5D",
x"4E28",
x"4DF2",
x"4DBC",
x"4D86",
x"4D50",
x"4D19",
x"4CE2",
x"4CAB",
x"4C73",
x"4C3B",
x"4C03",
x"4BCB",
x"4B92",
x"4B5A",
x"4B21",
x"4AE8",
x"4AAE",
x"4A75",
x"4A3B",
x"4A01",
x"49C7",
x"498D",
x"4953",
x"4918",
x"48DE",
x"48A3",
x"4868",
x"482D",
x"47F2",
x"47B7",
x"477C",
x"4740",
x"4705",
x"46CA",
x"468E",
x"4653",
x"4618",
x"45DC",
x"45A1",
x"4565",
x"452A",
x"44EE",
x"44B3",
x"4478",
x"443D",
x"4401",
x"43C6",
x"438B",
x"4350",
x"4315",
x"42DB",
x"42A0",
x"4265",
x"422B",
x"41F1",
x"41B6",
x"417C",
x"4143",
x"4109",
x"40CF",
x"4096",
x"405D",
x"4024",
x"3FEB",
x"3FB2",
x"3F7A",
x"3F41",
x"3F09",
x"3ED2",
x"3E9A",
x"3E63",
x"3E2B",
x"3DF4",
x"3DBE",
x"3D87",
x"3D51",
x"3D1B",
x"3CE5",
x"3CAF",
x"3C7A",
x"3C45",
x"3C10",
x"3BDB",
x"3BA7",
x"3B73",
x"3B3F",
x"3B0B",
x"3AD8",
x"3AA5",
x"3A72",
x"3A3F",
x"3A0D",
x"39DA",
x"39A8",
x"3977",
x"3945",
x"3914",
x"38E3",
x"38B2",
x"3881",
x"3851",
x"3821",
x"37F1",
x"37C1",
x"3791",
x"3762",
x"3733",
x"3704",
x"36D5",
x"36A6",
x"3678",
x"3649",
x"361B",
x"35ED",
x"35BF",
x"3592",
x"3564",
x"3537",
x"350A",
x"34DD",
x"34B0",
x"3483",
x"3456",
x"3429",
x"33FD",
x"33D0",
x"33A4",
x"3378",
x"334C",
x"3320",
x"32F4",
x"32C8",
x"329C",
x"3270",
x"3244",
x"3218",
x"31ED",
x"31C1",
x"3195",
x"316A",
x"313E",
x"3113",
x"30E7",
x"30BC",
x"3090",
x"3064",
x"3039",
x"300D",
x"2FE2",
x"2FB6",
x"2F8A",
x"2F5F",
x"2F33",
x"2F07",
x"2EDB",
x"2EAF",
x"2E83",
x"2E57",
x"2E2B",
x"2DFF",
x"2DD3",
x"2DA7",
x"2D7B",
x"2D4E",
x"2D22",
x"2CF5",
x"2CC9",
x"2C9C",
x"2C6F",
x"2C42",
x"2C15",
x"2BE8",
x"2BBB",
x"2B8E",
x"2B61",
x"2B33",
x"2B06",
x"2AD8",
x"2AAB",
x"2A7D",
x"2A4F",
x"2A21",
x"29F3",
x"29C5",
x"2997",
x"2968",
x"293A",
x"290B",
x"28DD",
x"28AE",
x"287F",
x"2850",
x"2821",
x"27F2",
x"27C3",
x"2794",
x"2764",
x"2735",
x"2706",
x"26D6",
x"26A6",
x"2676",
x"2647",
x"2617",
x"25E7",
x"25B7",
x"2586",
x"2556",
x"2526",
x"24F6",
x"24C5",
x"2495",
x"2464",
x"2433",
x"2403",
x"23D2",
x"23A1",
x"2370",
x"233F",
x"230E",
x"22DD",
x"22AC",
x"227B",
x"224A",
x"2218",
x"21E7",
x"21B6",
x"2184",
x"2153",
x"2121",
x"20EF",
x"20BE",
x"208C",
x"205A",
x"2028",
x"1FF7",
x"1FC5",
x"1F93",
x"1F61",
x"1F2F",
x"1EFD",
x"1ECA",
x"1E98",
x"1E66",
x"1E33",
x"1E01",
x"1DCF",
x"1D9C",
x"1D6A",
x"1D37",
x"1D04",
x"1CD1",
x"1C9F",
x"1C6C",
x"1C39",
x"1C06",
x"1BD3",
x"1B9F",
x"1B6C",
x"1B39",
x"1B05",
x"1AD2",
x"1A9E",
x"1A6A",
x"1A37",
x"1A03",
x"19CF",
x"199B",
x"1966",
x"1932",
x"18FE",
x"18C9",
x"1895",
x"1860",
x"182B",
x"17F6",
x"17C1",
x"178B",
x"1756",
x"1720",
x"16EB",
x"16B5",
x"167F",
x"1648",
x"1612",
x"15DC",
x"15A5",
x"156E",
x"1537",
x"1500",
x"14C9",
x"1491",
x"1459",
x"1421",
x"13E9",
x"13B1",
x"1379",
x"1340",
x"1307",
x"12CE",
x"1295",
x"125B",
x"1221",
x"11E8",
x"11AD",
x"1173",
x"1139",
x"10FE",
x"10C3",
x"1088",
x"104C",
x"1010",
x"0FD5",
x"0F98",
x"0F5C",
x"0F20",
x"0EE3",
x"0EA6",
x"0E69",
x"0E2B",
x"0DED",
x"0DAF",
x"0D71",
x"0D33",
x"0CF4",
x"0CB5",
x"0C76",
x"0C37",
x"0BF8",
x"0BB8",
x"0B78",
x"0B38",
x"0AF8",
x"0AB7",
x"0A76",
x"0A35",
x"09F4",
x"09B3",
x"0971",
x"092F",
x"08EE",
x"08AB",
x"0869",
x"0827",
x"07E4",
x"07A1",
x"075E",
x"071B",
x"06D8",
x"0694",
x"0651",
x"060D",
x"05C9",
x"0585",
x"0541",
x"04FD",
x"04B8",
x"0474",
x"042F",
x"03EB",
x"03A6",
x"0361",
x"031C",
x"02D7",
x"0292",
x"024D",
x"0208",
x"01C2",
x"017D",
x"0138",
x"00F2",
x"00AD",
x"0068",
x"0022",
x"FFDE",
x"FF98",
x"FF53",
x"FF0E",
x"FEC8",
x"FE83",
x"FE3E",
x"FDF8",
x"FDB3",
x"FD6E",
x"FD29",
x"FCE4",
x"FC9F",
x"FC5A",
x"FC15",
x"FBD1",
x"FB8C",
x"FB48",
x"FB03",
x"FABF",
x"FA7B",
x"FA37",
x"F9F3",
x"F9AF",
x"F96C",
x"F928",
x"F8E5",
x"F8A2",
x"F85F",
x"F81C",
x"F7D9",
x"F797",
x"F755",
x"F712",
x"F6D1",
x"F68F",
x"F64D",
x"F60C",
x"F5CB",
x"F58A",
x"F549",
x"F508",
x"F4C8",
x"F488",
x"F448",
x"F408",
x"F3C9",
x"F38A",
x"F34B",
x"F30C",
x"F2CD",
x"F28F",
x"F251",
x"F213",
x"F1D5",
x"F197",
x"F15A",
x"F11D",
x"F0E0",
x"F0A4",
x"F068",
x"F02B",
x"EFF0",
x"EFB4",
x"EF78",
x"EF3D",
x"EF02",
x"EEC7",
x"EE8D",
x"EE53",
x"EE18",
x"EDDF",
x"EDA5",
x"ED6B",
x"ED32",
x"ECF9",
x"ECC0",
x"EC87",
x"EC4F",
x"EC17",
x"EBDF",
x"EBA7",
x"EB6F",
x"EB37",
x"EB00",
x"EAC9",
x"EA92",
x"EA5B",
x"EA24",
x"E9EE",
x"E9B8",
x"E981",
x"E94B",
x"E915",
x"E8E0",
x"E8AA",
x"E875",
x"E83F",
x"E80A",
x"E7D5",
x"E7A0",
x"E76B",
x"E737",
x"E702",
x"E6CE",
x"E69A",
x"E665",
x"E631",
x"E5FD",
x"E5C9",
x"E596",
x"E562",
x"E52E",
x"E4FB",
x"E4C7",
x"E494",
x"E461",
x"E42D",
x"E3FA",
x"E3C7",
x"E394",
x"E361",
x"E32F",
x"E2FC",
x"E2C9",
x"E296",
x"E264",
x"E231",
x"E1FF",
x"E1CD",
x"E19A",
x"E168",
x"E136",
x"E103",
x"E0D1",
x"E09F",
x"E06D",
x"E03B",
x"E009",
x"DFD8",
x"DFA6",
x"DF74",
x"DF42",
x"DF11",
x"DEDF",
x"DEAD",
x"DE7C",
x"DE4A",
x"DE19",
x"DDE8",
x"DDB6",
x"DD85",
x"DD54",
x"DD23",
x"DCF2",
x"DCC1",
x"DC90",
x"DC5F",
x"DC2E",
x"DBFD",
x"DBCD",
x"DB9C",
x"DB6B",
x"DB3B",
x"DB0A",
x"DADA",
x"DAAA",
x"DA7A",
x"DA49",
x"DA19",
x"D9E9",
x"D9B9",
x"D98A",
x"D95A",
x"D92A",
x"D8FA",
x"D8CB",
x"D89C",
x"D86C",
x"D83D",
x"D80E",
x"D7DF",
x"D7B0",
x"D781",
x"D752",
x"D723",
x"D6F5",
x"D6C6",
x"D698",
x"D669",
x"D63B",
x"D60D",
x"D5DF",
x"D5B1",
x"D583",
x"D555",
x"D528",
x"D4FA",
x"D4CD",
x"D49F",
x"D472",
x"D445",
x"D418",
x"D3EB",
x"D3BE",
x"D391",
x"D364",
x"D337",
x"D30B",
x"D2DE",
x"D2B2",
x"D285",
x"D259",
x"D22D",
x"D201",
x"D1D5",
x"D1A9",
x"D17D",
x"D151",
x"D125",
x"D0F9",
x"D0CD",
x"D0A1",
x"D076",
x"D04A",
x"D01E",
x"CFF3",
x"CFC7",
x"CF9C",
x"CF70",
x"CF44",
x"CF19",
x"CEED",
x"CEC2",
x"CE96",
x"CE6B",
x"CE3F",
x"CE13",
x"CDE8",
x"CDBC",
x"CD90",
x"CD64",
x"CD38",
x"CD0C",
x"CCE0",
x"CCB4",
x"CC88",
x"CC5C",
x"CC30",
x"CC03",
x"CBD7",
x"CBAA",
x"CB7D",
x"CB50",
x"CB23",
x"CAF6",
x"CAC9",
x"CA9C",
x"CA6E",
x"CA41",
x"CA13",
x"C9E5",
x"C9B7",
x"C988",
x"C95A",
x"C92B",
x"C8FC",
x"C8CD",
x"C89E",
x"C86F",
x"C83F",
x"C80F",
x"C7DF",
x"C7AF",
x"C77F",
x"C74E",
x"C71D",
x"C6EC",
x"C6BB",
x"C689",
x"C658",
x"C626",
x"C5F3",
x"C5C1",
x"C58E",
x"C55B",
x"C528",
x"C4F5",
x"C4C1",
x"C48D",
x"C459",
x"C425",
x"C3F0",
x"C3BB",
x"C386",
x"C351",
x"C31B",
x"C2E5",
x"C2AF",
x"C279",
x"C242",
x"C20C",
x"C1D5",
x"C19D",
x"C166",
x"C12E",
x"C0F7",
x"C0BF",
x"C086",
x"C04E",
x"C015",
x"BFDC",
x"BFA3",
x"BF6A",
x"BF31",
x"BEF7",
x"BEBD",
x"BE84",
x"BE4A",
x"BE0F",
x"BDD5",
x"BD9B",
x"BD60",
x"BD25",
x"BCEB",
x"BCB0",
x"BC75",
x"BC3A",
x"BBFF",
x"BBC3",
x"BB88",
x"BB4D",
x"BB12",
x"BAD6",
x"BA9B",
x"BA5F",
x"BA24",
x"B9E8",
x"B9AD",
x"B972",
x"B936",
x"B8FB",
x"B8C0",
x"B884",
x"B849",
x"B80E",
x"B7D3",
x"B798",
x"B75D",
x"B722",
x"B6E8",
x"B6AD",
x"B673",
x"B639",
x"B5FF",
x"B5C5",
x"B58B",
x"B552",
x"B518",
x"B4DF",
x"B4A6",
x"B46E",
x"B435",
x"B3FD",
x"B3C5",
x"B38D",
x"B355",
x"B31E",
x"B2E7",
x"B2B0",
x"B27A",
x"B244",
x"B20E",
x"B1D8",
x"B1A3",
x"B16E",
x"B139",
x"B105",
x"B0D1",
x"B09D",
x"B069",
x"B036",
x"B004",
x"AFD1",
x"AF9F",
x"AF6D",
x"AF3C",
x"AF0B",
x"AEDA",
x"AEAA",
x"AE79",
x"AE4A",
x"AE1A",
x"ADEB",
x"ADBD",
x"AD8E",
x"AD60",
x"AD33",
x"AD05",
x"ACD8",
x"ACAC",
x"AC80",
x"AC54",
x"AC28",
x"ABFD",
x"ABD2",
x"ABA7",
x"AB7C",
x"AB52",
x"AB29",
x"AAFF",
x"AAD6",
x"AAAD",
x"AA84",
x"AA5C",
x"AA34",
x"AA0C",
x"A9E4",
x"A9BD",
x"A996",
x"A96F",
x"A948",
x"A921",
x"A8FB",
x"A8D5",
x"A8AF",
x"A889",
x"A864",
x"A83E",
x"A819",
x"A7F4",
x"A7CF",
x"A7AA",
x"A785",
x"A760",
x"A73C",
x"A717",
x"A6F3",
x"A6CE",
x"A6AA",
x"A686",
x"A661",
x"A63D",
x"A619",
x"A5F5",
x"A5D0",
x"A5AC",
x"A588",
x"A563",
x"A53F",
x"A51A",
x"A4F6",
x"A4D1",
x"A4AC",
x"A488",
x"A463",
x"A43E",
x"A418",
x"A3F3",
x"A3CE",
x"A3A8",
x"A382",
x"A35C",
x"A336",
x"A310",
x"A2E9",
x"A2C2",
x"A29C",
x"A274",
x"A24D",
x"A226",
x"A1FE",
x"A1D6",
x"A1AD",
x"A185",
x"A15C",
x"A133",
x"A10A",
x"A0E0",
x"A0B7",
x"A08D",
x"A062",
x"A038",
x"A00D",
x"9FE2",
x"9FB6",
x"9F8A",
x"9F5E",
x"9F32",
x"9F06",
x"9ED9",
x"9EAC",
x"9E7E",
x"9E51",
x"9E23",
x"9DF5",
x"9DC6",
x"9D97",
x"9D68",
x"9D39",
x"9D09",
x"9CDA",
x"9CAA",
x"9C79",
x"9C49",
x"9C18",
x"9BE7",
x"9BB6",
x"9B84",
x"9B52",
x"9B20",
x"9AEE",
x"9ABC",
x"9A89",
x"9A57",
x"9A24",
x"99F1",
x"99BE",
x"998A",
x"9957",
x"9923",
x"98EF",
x"98BB",
x"9887",
x"9853",
x"981E",
x"97EA",
x"97B5",
x"9781",
x"974C",
x"9718",
x"96E3",
x"96AE",
x"9679",
x"9644",
x"960F",
x"95DA",
x"95A6",
x"9571",
x"953C",
x"9507",
x"94D2",
x"949D",
x"9469",
x"9434",
x"93FF",
x"93CB",
x"9396",
x"9362",
x"932D",
x"92F9",
x"92C5",
x"9291",
x"925D",
x"922A",
x"91F6",
x"91C3",
x"918F",
x"915C",
x"9129",
x"90F6",
x"90C4",
x"9091",
x"905F",
x"902D",
x"8FFB",
x"8FC9",
x"8F97",
x"8F66",
x"8F35",
x"8F04",
x"8ED3",
x"8EA2",
x"8E72",
x"8E41",
x"8E11",
x"8DE2",
x"8DB2",
x"8D83",
x"8D53",
x"8D24",
x"8CF5",
x"8CC7",
x"8C98",
x"8C6A",
x"8C3C",
x"8C0E",
x"8BE1",
x"8BB3",
x"8B86",
x"8B59",
x"8B2C",
x"8AFF",
x"8AD2",
x"8AA6",
x"8A79",
x"8A4D",
x"8A21",
x"89F5",
x"89CA",
x"899E",
x"8972",
x"8947",
x"891C",
x"88F0",
x"88C5",
x"889A",
x"886F",
x"8844",
x"881A",
x"87EF",
x"87C4",
x"8799",
x"876F",
x"8744",
x"8719",
x"86EF",
x"86C4",
x"869A",
x"866F",
x"8644",
x"861A",
x"85EF",
x"85C4",
x"8599",
x"856F",
x"8544",
x"8519",
x"84ED",
x"84C2",
x"8497",
x"846C",
x"8440",
x"8415",
x"83E9",
x"83BD",
x"8391",
x"8365",
x"8339",
x"830C",
x"82E0",
x"82B3",
x"8286",
x"8259",
x"822C",
x"81FE",
x"81D1",
x"81A3",
x"8175",
x"8147",
x"8119",
x"80EA",
x"80BB",
x"808D",
x"805E",
x"802E",
x"7FFF",
x"7FCF",
x"7F9F",
x"7F6F",
x"7F3F",
x"7F0F",
x"7EDE",
x"7EAD",
x"7E7C",
x"7E4B",
x"7E1A",
x"7DE9",
x"7DB7",
x"7D85",
x"7D53",
x"7D21",
x"7CEF",
x"7CBD",
x"7C8A",
x"7C58",
x"7C25",
x"7BF2",
x"7BBF",
x"7B8C",
x"7B59",
x"7B26",
x"7AF2",
x"7ABF",
x"7A8C",
x"7A58",
x"7A25",
x"79F1",
x"79BE",
x"798A",
x"7957",
x"7923",
x"78F0",
x"78BC",
x"7889",
x"7856",
x"7822",
x"77EF",
x"77BC",
x"7789",
x"7756",
x"7723",
x"76F0",
x"76BE",
x"768B",
x"7659",
x"7627",
x"75F5",
x"75C3",
x"7592",
x"7561",
x"7530",
x"74FF",
x"74CE",
x"749E",
x"746D",
x"743D",
x"740E",
x"73DE",
x"73AF",
x"7380",
x"7352",
x"7324",
x"72F6",
x"72C8",
x"729B",
x"726E",
x"7241",
x"7215",
x"71E9",
x"71BD",
x"7192",
x"7167",
x"713C",
x"7111",
x"70E7",
x"70BE",
x"7094",
x"706B",
x"7042",
x"701A",
x"6FF2",
x"6FCA",
x"6FA2",
x"6F7B",
x"6F54",
x"6F2D",
x"6F07",
x"6EE1",
x"6EBB",
x"6E96",
x"6E70",
x"6E4B",
x"6E26",
x"6E02",
x"6DDD",
x"6DB9",
x"6D95",
x"6D71",
x"6D4D",
x"6D29",
x"6D06",
x"6CE2",
x"6CBF",
x"6C9B",
x"6C78",
x"6C55",
x"6C32",
x"6C0E",
x"6BEB",
x"6BC8",
x"6BA4",
x"6B81",
x"6B5D",
x"6B39",
x"6B16",
x"6AF2",
x"6ACD",
x"6AA9",
x"6A84",
x"6A5F",
x"6A3A",
x"6A15",
x"69EF",
x"69C8",
x"69A2",
x"697B",
x"6954",
x"692C",
x"6904",
x"68DB",
x"68B2",
x"6888",
x"685E",
x"6833",
x"6807",
x"67DB",
x"67AF",
x"6781",
x"6753",
x"6725",
x"66F5",
x"66C5",
x"6694",
x"6663",
x"6631",
x"65FE",
x"65CA",
x"6595",
x"655F",
x"6529",
x"64F2",
x"64BA",
x"6481",
x"6447",
x"640D",
x"63D1",
x"6395",
x"6358",
x"631A",
x"62DB",
x"629B",
x"625A",
x"6219",
x"61D6",
x"6193",
x"614F",
x"6109",
x"60C4",
x"607D",
x"6035",
x"5FED",
x"5FA4",
x"5F5A",
x"5F0F",
x"5EC4",
x"5E78",
x"5E2B",
x"5DDE",
x"5D90",
x"5D41",
x"5CF2",
x"5CA3",
x"5C52",
x"5C02",
x"5BB1",
x"5B5F",
x"5B0E",
x"5ABC",
x"5A69",
x"5A17",
x"59C4",
x"5971",
x"591F",
x"58CC",
x"5879",
x"5826",
x"57D4",
x"5782",
x"5730",
x"56DE",
x"568D",
x"563D",
x"55ED",
x"559D",
x"554E",
x"5500",
x"54B3",
x"5467",
x"541C",
x"53D2",
x"5389",
x"5341",
x"52FB",
x"52B6",
x"5273",
x"5231",
x"51F1",
x"51B2",
x"5176",
x"513B",
x"5103",
x"50CD",
x"5098",
x"5067",
x"5037",
x"500A",
x"4FE0",
x"4FB9",
x"4F94",
x"4F72",
x"4F53",
x"4F38",
x"4F1F",
x"4F0A",
x"4EF8",
x"4EEA",
x"4EE0",
x"4ED9",
x"4ED6",
x"4ED6",
x"4EDB",
x"4EE4",
x"4EF1",
x"4F03",
x"4F19",
x"4F33",
x"4F52",
x"4F76",
x"4F9E",
x"4FCC",
x"4FFE",
x"5036",
x"5072",
x"50B4",
x"50FC",
x"5149",
x"519B",
x"51F3",
x"5250",
x"52B4",
x"531D",
x"538C",
x"5402",
x"547D",
x"54FF",
x"5587",
x"5615",
x"56A9",
x"5744",
x"57E6",
x"588E",
x"593D",
x"59F2",
x"5AAF",
x"5B72",
x"5C3C",
x"5D0D",
x"5DE5",
x"5EC3",
x"5FA9",
x"6096",
x"618A",
x"6286",
x"6388",
x"6492",
x"65A3",
x"66BB",
x"67DA",
x"6901",
x"6A2F",
x"6B64",
x"6CA0",
x"6DE4",
x"6F2F",
x"7082",
x"71DB",
x"733C",
x"74A4",
x"7614",
x"778B",
x"7908",
x"7A8E",
x"7C1A",
x"7DAD",
x"7F47",
x"80E9",
x"8291",
x"8440",
x"85F6",
x"87B3",
x"8977",
x"8B41",
x"8D12",
x"8EEA",
x"90C8",
x"92AC",
x"9497",
x"9688",
x"987F",
x"9A7C",
x"9C80",
x"9E89",
x"A098",
x"A2AD",
x"A4C7",
x"A6E7",
x"A90C",
x"AB37",
x"AD66",
x"AF9B",
x"B1D5",
x"B413",
x"B656",
x"B89E",
x"BAEA",
x"BD3B",
x"BF8F",
x"C1E8",
x"C444",
x"C6A5",
x"C909",
x"CB70",
x"CDDB",
x"D049",
x"D2BA",
x"D52E",
x"D7A4",
x"DA1D",
x"DC99",
x"DF17",
x"E197",
x"E419",
x"E69C",
x"E922",
x"EBA8",
x"EE31",
x"F0BA",
x"F344",
x"F5CF",
x"F85B",
x"FAE7",
x"FD74",
x"0000"

    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            dout <= lut(to_integer(unsigned(addr)));
        end if;
    end process;
end arch;
