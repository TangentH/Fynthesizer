Library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;
use IEEE.NUMERIC_STD.ALL; 

entity sine_lut is
    generic (
        DEPTH : integer := 2048;  -- ���ñ�����ȣ��ɴ�?2048������
        WIDTH : integer := 16     -- ÿ������16λ��
    );
    port (
        clk   : in  std_logic;
        addr  : in  std_logic_vector(10 downto 0); -- 2048����������ַΪ11λ��
        dout  : out std_logic_vector(WIDTH-1 downto 0)
    );
end sine_lut;

architecture arch of sine_lut is
    type lut_array is array(0 to DEPTH-1) of std_logic_vector(WIDTH-1 downto 0);
    signal lut: lut_array := (
    x"4000", x"4032", x"4064", x"4096", x"40C9", x"40FB", x"412D", x"415F", x"4192", x"41C4", x"41F6", x"4228", x"425B", x"428D", x"42BF", x"42F1", x"4323", x"4356", x"4388", x"43BA", x"43EC", x"441E", x"4451", x"4483", x"44B5", x"44E7", x"4519", x"454B", x"457D", x"45AF", x"45E1", x"4613", x"4645", x"4677", x"46A9", x"46DB", x"470D", x"473F", x"4771", x"47A3", x"47D5", x"4807", x"4839", x"486B", x"489C", x"48CE", x"4900", x"4932", x"4964", x"4995", x"49C7", x"49F9", x"4A2A", x"4A5C", x"4A8D", x"4ABF", x"4AF1", x"4B22", x"4B54", x"4B85", x"4BB6", x"4BE8", x"4C19", x"4C4B", x"4C7C", x"4CAD", x"4CDE", x"4D10", x"4D41", x"4D72", x"4DA3", x"4DD4", x"4E05", x"4E36", x"4E67", x"4E98", x"4EC9", x"4EFA", x"4F2B", x"4F5C", x"4F8C", x"4FBD", x"4FEE", x"501F", x"504F", x"5080", x"50B0", x"50E1", x"5111", x"5142", x"5172", x"51A2", x"51D3", x"5203", x"5233", x"5263", x"5294", x"52C4", x"52F4", x"5324", x"5354", x"5383", x"53B3", x"53E3", x"5413", x"5443", x"5472", x"54A2", x"54D1", x"5501", x"5530", x"5560", x"558F", x"55BE", x"55EE", x"561D", x"564C", x"567B", x"56AA", x"56D9", x"5708", x"5737", x"5766", x"5794", x"57C3", x"57F2", x"5820", x"584F", x"587D", x"58AC", x"58DA", x"5908", x"5937", x"5965", x"5993", x"59C1", x"59EF", x"5A1D", x"5A4B", x"5A79", x"5AA6", x"5AD4", x"5B02", x"5B2F", x"5B5D", x"5B8A", x"5BB7", x"5BE5", x"5C12", x"5C3F", x"5C6C", x"5C99", x"5CC6", x"5CF3", x"5D20", x"5D4C", x"5D79", x"5DA6", x"5DD2", x"5DFE", x"5E2B", x"5E57", x"5E83", x"5EB0", x"5EDC", x"5F08", x"5F34", x"5F5F", x"5F8B", x"5FB7", x"5FE2", x"600E", x"6039", x"6065", x"6090", x"60BB", x"60E7", x"6112", x"613D", x"6168", x"6192", x"61BD", x"61E8", x"6212", x"623D", x"6267", x"6292", x"62BC", x"62E6", x"6310", x"633A", x"6364", x"638E", x"63B8", x"63E1", x"640B", x"6434", x"645E", x"6487", x"64B0", x"64DA", x"6503", x"652C", x"6554", x"657D", x"65A6", x"65CF", x"65F7", x"661F", x"6648", x"6670", x"6698", x"66C0", x"66E8", x"6710", x"6738", x"675F", x"6787", x"67AF", x"67D6", x"67FD", x"6824", x"684B", x"6872", x"6899", x"68C0", x"68E7", x"690E", x"6934", x"695A", x"6981", x"69A7", x"69CD", x"69F3", x"6A19", x"6A3F", x"6A65", x"6A8A", x"6AB0", x"6AD5", x"6AFA", x"6B20", x"6B45", x"6B6A", x"6B8E", x"6BB3", x"6BD8", x"6BFC", x"6C21", x"6C45", x"6C6A", x"6C8E", x"6CB2", x"6CD6", x"6CF9", x"6D1D", x"6D41", x"6D64", x"6D88", x"6DAB", x"6DCE", x"6DF1", x"6E14", x"6E37", x"6E5A", x"6E7C", x"6E9F", x"6EC1", x"6EE3", x"6F05", x"6F28", x"6F49", x"6F6B", x"6F8D", x"6FAF", x"6FD0", x"6FF1", x"7013", x"7034", x"7055", x"7076", x"7096", x"70B7", x"70D8", x"70F8", x"7118", x"7138", x"7159", x"7179", x"7198", x"71B8", x"71D8", x"71F7", x"7216", x"7236", x"7255", x"7274", x"7293", x"72B1", x"72D0", x"72EE", x"730D", x"732B", x"7349", x"7367", x"7385", x"73A3", x"73C1", x"73DE", x"73FB", x"7419", x"7436", x"7453", x"7470", x"748C", x"74A9", x"74C6", x"74E2", x"74FE", x"751A", x"7536", x"7552", x"756E", x"7589", x"75A5", x"75C0", x"75DC", x"75F7", x"7612", x"762C", x"7647", x"7662", x"767C", x"7696", x"76B1", x"76CB", x"76E5", x"76FE", x"7718", x"7731", x"774B", x"7764", x"777D", x"7796", x"77AF", x"77C8", x"77E0", x"77F9", x"7811", x"7829", x"7841", x"7859", x"7871", x"7889", x"78A0", x"78B7", x"78CF", x"78E6", x"78FD", x"7913", x"792A", x"7941", x"7957", x"796D", x"7983", x"7999", x"79AF", x"79C5", x"79DA", x"79F0", x"7A05", x"7A1A", x"7A2F", x"7A44", x"7A59", x"7A6D", x"7A82", x"7A96", x"7AAA", x"7ABE", x"7AD2", x"7AE6", x"7AFA", x"7B0D", x"7B20", x"7B34", x"7B47", x"7B59", x"7B6C", x"7B7F", x"7B91", x"7BA3", x"7BB6", x"7BC8", x"7BDA", x"7BEB", x"7BFD", x"7C0E", x"7C20", x"7C31", x"7C42", x"7C53", x"7C63", x"7C74", x"7C84", x"7C95", x"7CA5", x"7CB5", x"7CC5", x"7CD4", x"7CE4", x"7CF3", x"7D02", x"7D12", x"7D21", x"7D2F", x"7D3E", x"7D4D", x"7D5B", x"7D69", x"7D77", x"7D85", x"7D93", x"7DA1", x"7DAE", x"7DBB", x"7DC9", x"7DD6", x"7DE2", x"7DEF", x"7DFC", x"7E08", x"7E14", x"7E21", x"7E2D", x"7E38", x"7E44", x"7E50", x"7E5B", x"7E66", x"7E71", x"7E7C", x"7E87", x"7E92", x"7E9C", x"7EA7", x"7EB1", x"7EBB", x"7EC5", x"7ECE", x"7ED8", x"7EE1", x"7EEB", x"7EF4", x"7EFD", x"7F06", x"7F0E", x"7F17", x"7F1F", x"7F27", x"7F2F", x"7F37", x"7F3F", x"7F47", x"7F4E", x"7F55", x"7F5D", x"7F64", x"7F6A", x"7F71", x"7F78", x"7F7E", x"7F84", x"7F8A", x"7F90", x"7F96", x"7F9C", x"7FA1", x"7FA6", x"7FAC", x"7FB1", x"7FB5", x"7FBA", x"7FBF", x"7FC3", x"7FC7", x"7FCB", x"7FCF", x"7FD3", x"7FD7", x"7FDA", x"7FDE", x"7FE1", x"7FE4", x"7FE7", x"7FE9", x"7FEC", x"7FEE", x"7FF0", x"7FF2", x"7FF4", x"7FF6", x"7FF8", x"7FF9", x"7FFB", x"7FFC", x"7FFD", x"7FFE", x"7FFE", x"7FFF", x"7FFF", x"7FFF", x"8000", x"7FFF", x"7FFF", x"7FFF", x"7FFE", x"7FFE", x"7FFD", x"7FFC", x"7FFB", x"7FF9", x"7FF8", x"7FF6", x"7FF4", x"7FF2", x"7FF0", x"7FEE", x"7FEC", x"7FE9", x"7FE7", x"7FE4", x"7FE1", x"7FDE", x"7FDA", x"7FD7", x"7FD3", x"7FCF", x"7FCB", x"7FC7", x"7FC3", x"7FBF", x"7FBA", x"7FB5", x"7FB1", x"7FAC", x"7FA6", x"7FA1", x"7F9C", x"7F96", x"7F90", x"7F8A", x"7F84", x"7F7E", x"7F78", x"7F71", x"7F6A", x"7F64", x"7F5D", x"7F55", x"7F4E", x"7F47", x"7F3F", x"7F37", x"7F2F", x"7F27", x"7F1F", x"7F17", x"7F0E", x"7F06", x"7EFD", x"7EF4", x"7EEB", x"7EE1", x"7ED8", x"7ECE", x"7EC5", x"7EBB", x"7EB1", x"7EA7", x"7E9C", x"7E92", x"7E87", x"7E7C", x"7E71", x"7E66", x"7E5B", x"7E50", x"7E44", x"7E38", x"7E2D", x"7E21", x"7E14", x"7E08", x"7DFC", x"7DEF", x"7DE2", x"7DD6", x"7DC9", x"7DBB", x"7DAE", x"7DA1", x"7D93", x"7D85", x"7D77", x"7D69", x"7D5B", x"7D4D", x"7D3E", x"7D2F", x"7D21", x"7D12", x"7D02", x"7CF3", x"7CE4", x"7CD4", x"7CC5", x"7CB5", x"7CA5", x"7C95", x"7C84", x"7C74", x"7C63", x"7C53", x"7C42", x"7C31", x"7C20", x"7C0E", x"7BFD", x"7BEB", x"7BDA", x"7BC8", x"7BB6", x"7BA3", x"7B91", x"7B7F", x"7B6C", x"7B59", x"7B47", x"7B34", x"7B20", x"7B0D", x"7AFA", x"7AE6", x"7AD2", x"7ABE", x"7AAA", x"7A96", x"7A82", x"7A6D", x"7A59", x"7A44", x"7A2F", x"7A1A", x"7A05", x"79F0", x"79DA", x"79C5", x"79AF", x"7999", x"7983", x"796D", x"7957", x"7941", x"792A", x"7913", x"78FD", x"78E6", x"78CF", x"78B7", x"78A0", x"7889", x"7871", x"7859", x"7841", x"7829", x"7811", x"77F9", x"77E0", x"77C8", x"77AF", x"7796", x"777D", x"7764", x"774B", x"7731", x"7718", x"76FE", x"76E5", x"76CB", x"76B1", x"7696", x"767C", x"7662", x"7647", x"762C", x"7612", x"75F7", x"75DC", x"75C0", x"75A5", x"7589", x"756E", x"7552", x"7536", x"751A", x"74FE", x"74E2", x"74C6", x"74A9", x"748C", x"7470", x"7453", x"7436", x"7419", x"73FB", x"73DE", x"73C1", x"73A3", x"7385", x"7367", x"7349", x"732B", x"730D", x"72EE", x"72D0", x"72B1", x"7293", x"7274", x"7255", x"7236", x"7216", x"71F7", x"71D8", x"71B8", x"7198", x"7179", x"7159", x"7138", x"7118", x"70F8", x"70D8", x"70B7", x"7096", x"7076", x"7055", x"7034", x"7013", x"6FF1", x"6FD0", x"6FAF", x"6F8D", x"6F6B", x"6F49", x"6F28", x"6F05", x"6EE3", x"6EC1", x"6E9F", x"6E7C", x"6E5A", x"6E37", x"6E14", x"6DF1", x"6DCE", x"6DAB", x"6D88", x"6D64", x"6D41", x"6D1D", x"6CF9", x"6CD6", x"6CB2", x"6C8E", x"6C6A", x"6C45", x"6C21", x"6BFC", x"6BD8", x"6BB3", x"6B8E", x"6B6A", x"6B45", x"6B20", x"6AFA", x"6AD5", x"6AB0", x"6A8A", x"6A65", x"6A3F", x"6A19", x"69F3", x"69CD", x"69A7", x"6981", x"695A", x"6934", x"690E", x"68E7", x"68C0", x"6899", x"6872", x"684B", x"6824", x"67FD", x"67D6", x"67AF", x"6787", x"675F", x"6738", x"6710", x"66E8", x"66C0", x"6698", x"6670", x"6648", x"661F", x"65F7", x"65CF", x"65A6", x"657D", x"6554", x"652C", x"6503", x"64DA", x"64B0", x"6487", x"645E", x"6434", x"640B", x"63E1", x"63B8", x"638E", x"6364", x"633A", x"6310", x"62E6", x"62BC", x"6292", x"6267", x"623D", x"6212", x"61E8", x"61BD", x"6192", x"6168", x"613D", x"6112", x"60E7", x"60BB", x"6090", x"6065", x"6039", x"600E", x"5FE2", x"5FB7", x"5F8B", x"5F5F", x"5F34", x"5F08", x"5EDC", x"5EB0", x"5E83", x"5E57", x"5E2B", x"5DFE", x"5DD2", x"5DA6", x"5D79", x"5D4C", x"5D20", x"5CF3", x"5CC6", x"5C99", x"5C6C", x"5C3F", x"5C12", x"5BE5", x"5BB7", x"5B8A", x"5B5D", x"5B2F", x"5B02", x"5AD4", x"5AA6", x"5A79", x"5A4B", x"5A1D", x"59EF", x"59C1", x"5993", x"5965", x"5937", x"5908", x"58DA", x"58AC", x"587D", x"584F", x"5820", x"57F2", x"57C3", x"5794", x"5766", x"5737", x"5708", x"56D9", x"56AA", x"567B", x"564C", x"561D", x"55EE", x"55BE", x"558F", x"5560", x"5530", x"5501", x"54D1", x"54A2", x"5472", x"5443", x"5413", x"53E3", x"53B3", x"5383", x"5354", x"5324", x"52F4", x"52C4", x"5294", x"5263", x"5233", x"5203", x"51D3", x"51A2", x"5172", x"5142", x"5111", x"50E1", x"50B0", x"5080", x"504F", x"501F", x"4FEE", x"4FBD", x"4F8C", x"4F5C", x"4F2B", x"4EFA", x"4EC9", x"4E98", x"4E67", x"4E36", x"4E05", x"4DD4", x"4DA3", x"4D72", x"4D41", x"4D10", x"4CDE", x"4CAD", x"4C7C", x"4C4B", x"4C19", x"4BE8", x"4BB6", x"4B85", x"4B54", x"4B22", x"4AF1", x"4ABF", x"4A8D", x"4A5C", x"4A2A", x"49F9", x"49C7", x"4995", x"4964", x"4932", x"4900", x"48CE", x"489C", x"486B", x"4839", x"4807", x"47D5", x"47A3", x"4771", x"473F", x"470D", x"46DB", x"46A9", x"4677", x"4645", x"4613", x"45E1", x"45AF", x"457D", x"454B", x"4519", x"44E7", x"44B5", x"4483", x"4451", x"441E", x"43EC", x"43BA", x"4388", x"4356", x"4323", x"42F1", x"42BF", x"428D", x"425B", x"4228", x"41F6", x"41C4", x"4192", x"415F", x"412D", x"40FB", x"40C9", x"4096", x"4064", x"4032", x"4000", x"3FCD", x"3F9B", x"3F69", x"3F36", x"3F04", x"3ED2", x"3EA0", x"3E6D", x"3E3B", x"3E09", x"3DD7", x"3DA4", x"3D72", x"3D40", x"3D0E", x"3CDC", x"3CA9", x"3C77", x"3C45", x"3C13", x"3BE1", x"3BAE", x"3B7C", x"3B4A", x"3B18", x"3AE6", x"3AB4", x"3A82", x"3A50", x"3A1E", x"39EC", x"39BA", x"3988", x"3956", x"3924", x"38F2", x"38C0", x"388E", x"385C", x"382A", x"37F8", x"37C6", x"3794", x"3763", x"3731", x"36FF", x"36CD", x"369B", x"366A", x"3638", x"3606", x"35D5", x"35A3", x"3572", x"3540", x"350E", x"34DD", x"34AB", x"347A", x"3449", x"3417", x"33E6", x"33B4", x"3383", x"3352", x"3321", x"32EF", x"32BE", x"328D", x"325C", x"322B", x"31FA", x"31C9", x"3198", x"3167", x"3136", x"3105", x"30D4", x"30A3", x"3073", x"3042", x"3011", x"2FE0", x"2FB0", x"2F7F", x"2F4F", x"2F1E", x"2EEE", x"2EBD", x"2E8D", x"2E5D", x"2E2C", x"2DFC", x"2DCC", x"2D9C", x"2D6B", x"2D3B", x"2D0B", x"2CDB", x"2CAB", x"2C7C", x"2C4C", x"2C1C", x"2BEC", x"2BBC", x"2B8D", x"2B5D", x"2B2E", x"2AFE", x"2ACF", x"2A9F", x"2A70", x"2A41", x"2A11", x"29E2", x"29B3", x"2984", x"2955", x"2926", x"28F7", x"28C8", x"2899", x"286B", x"283C", x"280D", x"27DF", x"27B0", x"2782", x"2753", x"2725", x"26F7", x"26C8", x"269A", x"266C", x"263E", x"2610", x"25E2", x"25B4", x"2586", x"2559", x"252B", x"24FD", x"24D0", x"24A2", x"2475", x"2448", x"241A", x"23ED", x"23C0", x"2393", x"2366", x"2339", x"230C", x"22DF", x"22B3", x"2286", x"2259", x"222D", x"2201", x"21D4", x"21A8", x"217C", x"214F", x"2123", x"20F7", x"20CB", x"20A0", x"2074", x"2048", x"201D", x"1FF1", x"1FC6", x"1F9A", x"1F6F", x"1F44", x"1F18", x"1EED", x"1EC2", x"1E97", x"1E6D", x"1E42", x"1E17", x"1DED", x"1DC2", x"1D98", x"1D6D", x"1D43", x"1D19", x"1CEF", x"1CC5", x"1C9B", x"1C71", x"1C47", x"1C1E", x"1BF4", x"1BCB", x"1BA1", x"1B78", x"1B4F", x"1B25", x"1AFC", x"1AD3", x"1AAB", x"1A82", x"1A59", x"1A30", x"1A08", x"19E0", x"19B7", x"198F", x"1967", x"193F", x"1917", x"18EF", x"18C7", x"18A0", x"1878", x"1850", x"1829", x"1802", x"17DB", x"17B4", x"178D", x"1766", x"173F", x"1718", x"16F1", x"16CB", x"16A5", x"167E", x"1658", x"1632", x"160C", x"15E6", x"15C0", x"159A", x"1575", x"154F", x"152A", x"1505", x"14DF", x"14BA", x"1495", x"1471", x"144C", x"1427", x"1403", x"13DE", x"13BA", x"1395", x"1371", x"134D", x"1329", x"1306", x"12E2", x"12BE", x"129B", x"1277", x"1254", x"1231", x"120E", x"11EB", x"11C8", x"11A5", x"1183", x"1160", x"113E", x"111C", x"10FA", x"10D7", x"10B6", x"1094", x"1072", x"1050", x"102F", x"100E", x"0FEC", x"0FCB", x"0FAA", x"0F89", x"0F69", x"0F48", x"0F27", x"0F07", x"0EE7", x"0EC7", x"0EA6", x"0E86", x"0E67", x"0E47", x"0E27", x"0E08", x"0DE9", x"0DC9", x"0DAA", x"0D8B", x"0D6C", x"0D4E", x"0D2F", x"0D11", x"0CF2", x"0CD4", x"0CB6", x"0C98", x"0C7A", x"0C5C", x"0C3E", x"0C21", x"0C04", x"0BE6", x"0BC9", x"0BAC", x"0B8F", x"0B73", x"0B56", x"0B39", x"0B1D", x"0B01", x"0AE5", x"0AC9", x"0AAD", x"0A91", x"0A76", x"0A5A", x"0A3F", x"0A23", x"0A08", x"09ED", x"09D3", x"09B8", x"099D", x"0983", x"0969", x"094E", x"0934", x"091A", x"0901", x"08E7", x"08CE", x"08B4", x"089B", x"0882", x"0869", x"0850", x"0837", x"081F", x"0806", x"07EE", x"07D6", x"07BE", x"07A6", x"078E", x"0776", x"075F", x"0748", x"0730", x"0719", x"0702", x"06EC", x"06D5", x"06BE", x"06A8", x"0692", x"067C", x"0666", x"0650", x"063A", x"0625", x"060F", x"05FA", x"05E5", x"05D0", x"05BB", x"05A6", x"0592", x"057D", x"0569", x"0555", x"0541", x"052D", x"0519", x"0505", x"04F2", x"04DF", x"04CB", x"04B8", x"04A6", x"0493", x"0480", x"046E", x"045C", x"0449", x"0437", x"0425", x"0414", x"0402", x"03F1", x"03DF", x"03CE", x"03BD", x"03AC", x"039C", x"038B", x"037B", x"036A", x"035A", x"034A", x"033A", x"032B", x"031B", x"030C", x"02FD", x"02ED", x"02DE", x"02D0", x"02C1", x"02B2", x"02A4", x"0296", x"0288", x"027A", x"026C", x"025E", x"0251", x"0244", x"0236", x"0229", x"021D", x"0210", x"0203", x"01F7", x"01EB", x"01DE", x"01D2", x"01C7", x"01BB", x"01AF", x"01A4", x"0199", x"018E", x"0183", x"0178", x"016D", x"0163", x"0158", x"014E", x"0144", x"013A", x"0131", x"0127", x"011E", x"0114", x"010B", x"0102", x"00F9", x"00F1", x"00E8", x"00E0", x"00D8", x"00D0", x"00C8", x"00C0", x"00B8", x"00B1", x"00AA", x"00A2", x"009B", x"0095", x"008E", x"0087", x"0081", x"007B", x"0075", x"006F", x"0069", x"0063", x"005E", x"0059", x"0053", x"004E", x"004A", x"0045", x"0040", x"003C", x"0038", x"0034", x"0030", x"002C", x"0028", x"0025", x"0021", x"001E", x"001B", x"0018", x"0016", x"0013", x"0011", x"000F", x"000D", x"000B", x"0009", x"0007", x"0006", x"0004", x"0003", x"0002", x"0001", x"0001", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0000", x"0001", x"0001", x"0002", x"0003", x"0004", x"0006", x"0007", x"0009", x"000B", x"000D", x"000F", x"0011", x"0013", x"0016", x"0018", x"001B", x"001E", x"0021", x"0025", x"0028", x"002C", x"0030", x"0034", x"0038", x"003C", x"0040", x"0045", x"004A", x"004E", x"0053", x"0059", x"005E", x"0063", x"0069", x"006F", x"0075", x"007B", x"0081", x"0087", x"008E", x"0095", x"009B", x"00A2", x"00AA", x"00B1", x"00B8", x"00C0", x"00C8", x"00D0", x"00D8", x"00E0", x"00E8", x"00F1", x"00F9", x"0102", x"010B", x"0114", x"011E", x"0127", x"0131", x"013A", x"0144", x"014E", x"0158", x"0163", x"016D", x"0178", x"0183", x"018E", x"0199", x"01A4", x"01AF", x"01BB", x"01C7", x"01D2", x"01DE", x"01EB", x"01F7", x"0203", x"0210", x"021D", x"0229", x"0236", x"0244", x"0251", x"025E", x"026C", x"027A", x"0288", x"0296", x"02A4", x"02B2", x"02C1", x"02D0", x"02DE", x"02ED", x"02FD", x"030C", x"031B", x"032B", x"033A", x"034A", x"035A", x"036A", x"037B", x"038B", x"039C", x"03AC", x"03BD", x"03CE", x"03DF", x"03F1", x"0402", x"0414", x"0425", x"0437", x"0449", x"045C", x"046E", x"0480", x"0493", x"04A6", x"04B8", x"04CB", x"04DF", x"04F2", x"0505", x"0519", x"052D", x"0541", x"0555", x"0569", x"057D", x"0592", x"05A6", x"05BB", x"05D0", x"05E5", x"05FA", x"060F", x"0625", x"063A", x"0650", x"0666", x"067C", x"0692", x"06A8", x"06BE", x"06D5", x"06EC", x"0702", x"0719", x"0730", x"0748", x"075F", x"0776", x"078E", x"07A6", x"07BE", x"07D6", x"07EE", x"0806", x"081F", x"0837", x"0850", x"0869", x"0882", x"089B", x"08B4", x"08CE", x"08E7", x"0901", x"091A", x"0934", x"094E", x"0969", x"0983", x"099D", x"09B8", x"09D3", x"09ED", x"0A08", x"0A23", x"0A3F", x"0A5A", x"0A76", x"0A91", x"0AAD", x"0AC9", x"0AE5", x"0B01", x"0B1D", x"0B39", x"0B56", x"0B73", x"0B8F", x"0BAC", x"0BC9", x"0BE6", x"0C04", x"0C21", x"0C3E", x"0C5C", x"0C7A", x"0C98", x"0CB6", x"0CD4", x"0CF2", x"0D11", x"0D2F", x"0D4E", x"0D6C", x"0D8B", x"0DAA", x"0DC9", x"0DE9", x"0E08", x"0E27", x"0E47", x"0E67", x"0E86", x"0EA6", x"0EC7", x"0EE7", x"0F07", x"0F27", x"0F48", x"0F69", x"0F89", x"0FAA", x"0FCB", x"0FEC", x"100E", x"102F", x"1050", x"1072", x"1094", x"10B6", x"10D7", x"10FA", x"111C", x"113E", x"1160", x"1183", x"11A5", x"11C8", x"11EB", x"120E", x"1231", x"1254", x"1277", x"129B", x"12BE", x"12E2", x"1306", x"1329", x"134D", x"1371", x"1395", x"13BA", x"13DE", x"1403", x"1427", x"144C", x"1471", x"1495", x"14BA", x"14DF", x"1505", x"152A", x"154F", x"1575", x"159A", x"15C0", x"15E6", x"160C", x"1632", x"1658", x"167E", x"16A5", x"16CB", x"16F1", x"1718", x"173F", x"1766", x"178D", x"17B4", x"17DB", x"1802", x"1829", x"1850", x"1878", x"18A0", x"18C7", x"18EF", x"1917", x"193F", x"1967", x"198F", x"19B7", x"19E0", x"1A08", x"1A30", x"1A59", x"1A82", x"1AAB", x"1AD3", x"1AFC", x"1B25", x"1B4F", x"1B78", x"1BA1", x"1BCB", x"1BF4", x"1C1E", x"1C47", x"1C71", x"1C9B", x"1CC5", x"1CEF", x"1D19", x"1D43", x"1D6D", x"1D98", x"1DC2", x"1DED", x"1E17", x"1E42", x"1E6D", x"1E97", x"1EC2", x"1EED", x"1F18", x"1F44", x"1F6F", x"1F9A", x"1FC6", x"1FF1", x"201D", x"2048", x"2074", x"20A0", x"20CB", x"20F7", x"2123", x"214F", x"217C", x"21A8", x"21D4", x"2201", x"222D", x"2259", x"2286", x"22B3", x"22DF", x"230C", x"2339", x"2366", x"2393", x"23C0", x"23ED", x"241A", x"2448", x"2475", x"24A2", x"24D0", x"24FD", x"252B", x"2559", x"2586", x"25B4", x"25E2", x"2610", x"263E", x"266C", x"269A", x"26C8", x"26F7", x"2725", x"2753", x"2782", x"27B0", x"27DF", x"280D", x"283C", x"286B", x"2899", x"28C8", x"28F7", x"2926", x"2955", x"2984", x"29B3", x"29E2", x"2A11", x"2A41", x"2A70", x"2A9F", x"2ACF", x"2AFE", x"2B2E", x"2B5D", x"2B8D", x"2BBC", x"2BEC", x"2C1C", x"2C4C", x"2C7C", x"2CAB", x"2CDB", x"2D0B", x"2D3B", x"2D6B", x"2D9C", x"2DCC", x"2DFC", x"2E2C", x"2E5D", x"2E8D", x"2EBD", x"2EEE", x"2F1E", x"2F4F", x"2F7F", x"2FB0", x"2FE0", x"3011", x"3042", x"3073", x"30A3", x"30D4", x"3105", x"3136", x"3167", x"3198", x"31C9", x"31FA", x"322B", x"325C", x"328D", x"32BE", x"32EF", x"3321", x"3352", x"3383", x"33B4", x"33E6", x"3417", x"3449", x"347A", x"34AB", x"34DD", x"350E", x"3540", x"3572", x"35A3", x"35D5", x"3606", x"3638", x"366A", x"369B", x"36CD", x"36FF", x"3731", x"3763", x"3794", x"37C6", x"37F8", x"382A", x"385C", x"388E", x"38C0", x"38F2", x"3924", x"3956", x"3988", x"39BA", x"39EC", x"3A1E", x"3A50", x"3A82", x"3AB4", x"3AE6", x"3B18", x"3B4A", x"3B7C", x"3BAE", x"3BE1", x"3C13", x"3C45", x"3C77", x"3CA9", x"3CDC", x"3D0E", x"3D40", x"3D72", x"3DA4", x"3DD7", x"3E09", x"3E3B", x"3E6D", x"3EA0", x"3ED2", x"3F04", x"3F36", x"3F69", x"3F9B", x"3FCD"
    );
begin
    process(clk)
    begin
        if rising_edge(clk) then
            dout <= lut(to_integer(unsigned(addr)));
        end if;
    end process;
end arch;